* Spice description of sum5b_cougar
* Spice driver version -1209512284
* Date ( dd/mm/yyyy hh:mm:ss ): 26/10/2020 at 21:06:13

* INTERF a[0] a[1] a[2] a[3] a[4] b[0] b[1] b[2] b[3] b[4] ci co so[0] so[1] 
* INTERF so[2] so[3] so[4] vdd vss 


.subckt sum5b_cougar 274 187 159 86 73 273 266 258 249 246 267 42 268 166 162 74 31 278 239 
* NET 9 = a3_x2_4_sig
* NET 14 = no3_x1_5_sig
* NET 15 = not_b[3]
* NET 16 = not_a[3]
* NET 20 = inv_x2_3_sig
* NET 24 = not_aux0
* NET 26 = a2_x2_sig
* NET 27 = not_a[4]
* NET 30 = no3_x1_7_sig
* NET 31 = so[4]
* NET 38 = ao2o22_x2_sig
* NET 42 = co
* NET 45 = no3_x1_sig
* NET 48 = no3_x1_8_sig
* NET 50 = inv_x2_sig
* NET 56 = not_aux25
* NET 59 = no4_x1_3_sig
* NET 60 = na3_x1_sig
* NET 61 = no2_x1_2_sig
* NET 62 = aux26
* NET 64 = aux1
* NET 73 = a[4]
* NET 74 = so[3]
* NET 75 = not_a[2]
* NET 78 = no3_x1_4_sig
* NET 79 = no2_x1_sig
* NET 83 = no3_x1_3_sig
* NET 85 = aux18
* NET 86 = a[3]
* NET 87 = a3_x2_2_sig
* NET 91 = aux3
* NET 93 = inv_x2_2_sig
* NET 94 = not_aux26
* NET 95 = no4_x1_sig
* NET 98 = no4_x1_4_sig
* NET 102 = not_aux8
* NET 103 = not_aux10
* NET 109 = no3_x1_6_sig
* NET 113 = na2_x1_sig
* NET 125 = no3_x1_2_sig
* NET 126 = nao22_x1_sig
* NET 132 = no4_x1_2_sig
* NET 134 = a3_x2_3_sig
* NET 135 = nao22_x1_2_sig
* NET 137 = no4_x1_5_sig
* NET 140 = not_aux27
* NET 141 = inv_x2_4_sig
* NET 145 = not_aux18
* NET 147 = a4_x2_sig
* NET 148 = not_ci
* NET 149 = not_a[0]
* NET 152 = aux23
* NET 155 = aux8
* NET 159 = a[2]
* NET 162 = so[2]
* NET 166 = so[1]
* NET 168 = not_aux30
* NET 169 = aux29
* NET 175 = oa2a22_x2_sig
* NET 176 = mbk_buf_aux5
* NET 177 = xr2_x1_3_sig
* NET 181 = not_aux24
* NET 182 = aux5
* NET 185 = xr2_x1_2_sig
* NET 187 = a[1]
* NET 189 = aux4
* NET 199 = a3_x2_sig
* NET 203 = not_aux33
* NET 209 = o3_x2_sig
* NET 211 = not_aux32
* NET 213 = mbk_buf_not_aux12
* NET 217 = not_aux12
* NET 218 = not_aux28
* NET 220 = not_aux31
* NET 225 = not_aux4
* NET 228 = not_a[1]
* NET 232 = not_aux9
* NET 234 = mbk_buf_not_aux9
* NET 237 = aux10
* NET 239 = vss
* NET 240 = oa2a22_x2_2_sig
* NET 244 = xr2_x1_4_sig
* NET 246 = b[4]
* NET 248 = not_aux15
* NET 249 = b[3]
* NET 251 = xr2_x1_5_sig
* NET 254 = aux12
* NET 256 = not_b[2]
* NET 257 = mbk_buf_aux12
* NET 258 = b[2]
* NET 259 = not_b[1]
* NET 260 = not_aux14
* NET 261 = aux15
* NET 262 = not_aux5
* NET 265 = not_aux6
* NET 266 = b[1]
* NET 267 = ci
* NET 268 = so[0]
* NET 271 = not_b[0]
* NET 273 = b[0]
* NET 274 = a[0]
* NET 277 = xr2_x1_sig
* NET 278 = vdd
Mtr_00532 270 267 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00531 278 277 272 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00530 268 270 269 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00529 269 277 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00528 269 272 268 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00527 278 267 269 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00526 275 274 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00525 278 273 276 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00524 277 275 279 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00523 279 273 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00522 279 276 277 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00521 278 274 279 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00520 271 273 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00519 259 266 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00518 264 262 263 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00517 278 271 264 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00516 265 263 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00515 261 260 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00514 278 265 261 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00513 257 255 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00512 278 254 255 278 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00511 242 251 241 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00510 242 266 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00509 278 244 242 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00508 241 259 242 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00507 240 241 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00506 243 258 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00505 278 261 247 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00504 244 243 245 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00503 245 261 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00502 245 247 244 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00501 278 258 245 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00500 256 258 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00499 248 261 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00498 250 258 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00497 278 257 253 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00496 251 250 252 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00495 252 257 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00494 252 253 251 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00493 278 258 252 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00492 260 226 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00491 278 225 226 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00490 226 228 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00489 234 233 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00488 278 232 233 278 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00487 217 254 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00486 197 234 235 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00485 278 271 197 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00484 237 235 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00483 220 222 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00482 278 225 222 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00481 222 265 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00480 196 262 229 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00479 278 228 196 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00478 232 229 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00477 278 232 195 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00476 254 225 195 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00475 195 271 254 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00474 194 258 219 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00473 278 266 194 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00472 218 219 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00471 278 259 192 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00470 192 248 191 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00469 191 256 210 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00468 209 210 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00467 278 209 211 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00466 193 213 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00465 211 256 193 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00464 278 204 203 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00463 190 199 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00462 190 248 204 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00461 204 256 190 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00460 278 217 202 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00459 199 202 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00458 278 259 202 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00457 202 256 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00456 213 214 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00455 278 217 214 278 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00454 189 188 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00453 278 267 188 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00452 188 274 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00451 225 189 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00450 181 180 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00449 278 260 180 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00448 180 271 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00447 228 187 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00446 262 182 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00445 183 187 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00444 278 189 184 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00443 185 183 186 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00442 186 189 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00441 186 184 185 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00440 278 187 186 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00439 171 187 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00438 278 176 172 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00437 177 171 173 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00436 173 176 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00435 173 172 177 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00434 278 187 173 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00433 179 177 178 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00432 179 271 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00431 278 185 179 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00430 178 273 179 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00429 175 178 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00428 176 174 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00427 278 182 174 278 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00426 168 187 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00425 278 258 168 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00424 170 258 169 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00423 278 187 170 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00422 160 159 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00421 278 240 161 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00420 162 160 163 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00419 163 240 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00418 163 161 162 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00417 278 159 163 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00416 164 266 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00415 278 175 167 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00414 166 164 165 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00413 165 175 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00412 165 167 166 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00411 278 266 165 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00410 149 274 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00409 278 148 152 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00408 152 149 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00407 152 228 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00406 278 267 155 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00405 155 274 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00404 155 187 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00403 147 146 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00402 146 237 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00401 278 256 146 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00400 146 145 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00399 278 155 146 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00398 278 259 115 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00397 117 181 116 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00396 116 256 137 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00395 115 140 117 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00394 141 152 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00393 278 181 118 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00392 120 141 119 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00391 119 256 132 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00390 118 145 120 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00389 113 152 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00388 278 137 113 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00387 278 169 131 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00386 134 131 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00385 278 220 131 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 131 145 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00383 278 259 126 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00382 105 125 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00381 126 147 105 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00380 278 266 135 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00379 110 134 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00378 135 132 110 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00377 278 140 108 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00376 107 220 109 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00375 108 168 107 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00374 278 168 106 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00373 104 145 125 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00372 106 220 104 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00371 103 237 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00370 148 267 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00369 145 85 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00368 93 91 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00367 278 103 92 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00366 97 102 96 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00365 96 218 95 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00364 92 91 97 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00363 182 149 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00362 278 148 182 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00361 102 155 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00360 278 94 100 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00359 99 102 101 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00358 101 103 98 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00357 100 218 99 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00356 278 84 89 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00355 89 88 85 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00354 89 86 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00353 85 249 89 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00352 278 86 88 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00351 84 249 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00350 278 159 81 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00349 82 211 83 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00348 81 85 82 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00347 278 93 90 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00346 87 90 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00345 278 169 90 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00344 90 220 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00343 278 203 77 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00342 76 145 78 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00341 77 75 76 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00340 80 83 79 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00339 278 78 80 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00338 278 135 74 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00337 74 126 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00336 74 79 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00335 71 246 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 278 73 72 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00333 56 71 53 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00332 53 73 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00331 53 72 56 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00330 278 246 53 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00329 278 69 91 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00328 51 50 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00327 51 246 69 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00326 69 73 51 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00325 278 159 47 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00324 46 211 48 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00323 47 94 46 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00322 94 62 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00321 278 220 60 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00320 60 62 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00319 60 169 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00318 62 63 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00317 278 64 63 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00316 63 56 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00315 49 98 61 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00314 278 48 49 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00313 278 159 44 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00312 43 211 45 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00311 44 91 43 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00310 278 45 40 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00309 39 38 41 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00308 41 87 42 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00307 40 95 39 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00306 75 159 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00305 278 60 31 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00304 31 61 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 278 59 31 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00302 31 113 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 278 203 29 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00300 28 140 30 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00299 29 75 28 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00298 26 25 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00297 278 24 25 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00296 25 27 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 27 73 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00294 20 246 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00293 21 20 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 23 24 22 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 278 27 23 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 22 26 21 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 38 22 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00288 18 56 19 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00287 278 24 18 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00286 140 19 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00285 50 64 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00284 16 86 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00283 24 17 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00282 278 15 17 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 17 16 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 64 86 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00279 278 249 64 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 278 56 8 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 9 8 278 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00276 278 15 8 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 8 16 278 278 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 15 249 278 278 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00273 278 14 7 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00272 12 9 13 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00271 13 30 59 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00270 7 109 12 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00269 278 56 11 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00268 10 16 14 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00267 11 15 10 278 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00266 272 277 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00265 239 267 270 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00264 230 270 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00263 268 272 230 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 231 267 268 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 239 277 231 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 276 273 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00259 239 274 275 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00258 238 275 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00257 277 276 238 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00256 236 274 277 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00255 239 273 236 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00254 239 273 271 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00253 239 266 259 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00252 265 263 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00251 263 271 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00250 239 262 263 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00249 239 260 223 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00248 223 265 261 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00247 239 255 257 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00246 255 254 239 239 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00245 206 251 241 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00244 239 259 206 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00243 205 266 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00242 241 244 205 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00241 239 241 240 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00240 247 261 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00239 239 258 243 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00238 208 243 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 244 247 208 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 207 258 244 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00235 239 261 207 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 239 258 256 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00233 239 261 248 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 253 257 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00231 239 258 250 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00230 216 250 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 251 253 216 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00228 215 258 251 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00227 239 257 215 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00226 226 228 227 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00225 239 226 260 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00224 227 225 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00223 239 233 234 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00222 233 232 239 239 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00221 239 254 217 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 237 235 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 235 271 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00218 239 234 235 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00217 222 265 221 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 239 222 220 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00215 221 225 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00214 232 229 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 229 228 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00212 239 262 229 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00211 239 225 224 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00210 224 271 254 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00209 254 232 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00208 218 219 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 219 266 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00206 239 258 219 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00205 210 256 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00204 210 259 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00203 239 248 210 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00202 239 210 209 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 212 213 211 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 211 256 212 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 212 209 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 203 204 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 239 199 204 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00196 200 248 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00195 204 256 200 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00194 239 202 199 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00193 198 217 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 201 256 198 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00191 202 259 201 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00190 239 214 213 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00189 214 217 239 239 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00188 188 274 158 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00187 239 188 189 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00186 158 267 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00185 239 189 225 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00184 180 271 144 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 239 180 181 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00182 144 260 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00181 239 187 228 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 239 182 262 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 184 189 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00178 239 187 183 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00177 154 183 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 185 184 154 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 153 187 185 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 239 189 153 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 172 176 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00172 239 187 171 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00171 139 171 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 177 172 139 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 138 187 177 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 239 176 138 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 143 177 178 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00166 239 273 143 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00165 142 271 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00164 178 185 142 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00163 239 178 175 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 239 174 176 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 174 182 239 239 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00160 239 187 136 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 136 258 168 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 169 187 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00157 239 258 169 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00156 161 240 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00155 239 159 160 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00154 124 160 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00153 162 161 124 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 128 159 162 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 239 240 128 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 167 175 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00149 239 266 164 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00148 130 164 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 166 167 130 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 129 266 166 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00145 239 175 129 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00144 239 274 149 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00143 239 228 151 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 151 148 150 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 150 149 152 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 239 187 156 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 156 267 157 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 157 274 155 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 122 145 121 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 239 237 123 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 121 155 146 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 123 256 122 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00133 239 146 147 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00132 137 259 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00131 239 256 137 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00130 239 140 137 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00129 137 181 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00128 239 152 141 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00127 132 181 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00126 239 256 132 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00125 239 145 132 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00124 132 141 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00123 239 152 114 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00122 114 137 113 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00121 239 131 134 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 112 169 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 111 145 112 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 131 220 111 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 127 125 126 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 126 147 127 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 127 259 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 133 134 135 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 135 132 133 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 133 266 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 239 168 109 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00110 109 140 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00109 109 220 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00108 239 220 125 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 125 168 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00106 125 145 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00105 239 237 103 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 239 267 148 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 239 85 145 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 239 91 93 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 95 103 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00100 239 218 95 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00099 239 91 95 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00098 95 102 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00097 239 149 70 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 70 148 182 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 239 155 102 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 98 94 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00093 239 103 98 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00092 239 218 98 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00091 98 102 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00090 239 86 66 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 66 84 85 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 85 88 65 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 65 249 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 239 249 84 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00085 88 86 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00084 239 85 83 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00083 83 159 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00082 83 211 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00081 239 90 87 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 68 93 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 67 220 68 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 90 169 67 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 239 75 78 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00076 78 203 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00075 78 145 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00074 79 78 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00073 239 83 79 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00072 239 79 58 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 58 135 57 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 57 126 74 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 72 73 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00068 239 246 71 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00067 55 71 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 56 72 55 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 54 246 56 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 239 73 54 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 91 69 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 239 50 69 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00061 52 246 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00060 69 73 52 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00059 239 94 48 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00058 48 159 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00057 48 211 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 239 62 94 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 239 169 36 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 36 220 35 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 35 62 60 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 63 56 37 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 239 63 62 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 37 64 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 61 48 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00048 239 98 61 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 239 91 45 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 45 159 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 45 211 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00044 42 45 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00043 239 87 42 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00042 239 95 42 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00041 42 38 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00040 239 159 75 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 239 113 34 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 34 60 32 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 32 61 33 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 33 59 31 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 239 75 30 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 30 203 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 30 140 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 25 27 6 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 239 25 26 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 6 24 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 239 73 27 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 239 246 20 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 5 24 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00026 239 27 5 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00025 5 20 22 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00024 22 26 5 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 239 22 38 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 140 19 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 19 24 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 239 56 19 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00019 239 64 50 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 239 86 16 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 17 16 4 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 239 17 24 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 4 15 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 239 86 3 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 3 249 64 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 239 8 9 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 1 56 239 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 2 16 1 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 8 15 2 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 239 249 15 239 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 59 14 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 239 30 59 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 239 109 59 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 59 9 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 239 15 14 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 14 56 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 14 16 239 239 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C281 5 239 7.43e-15
C277 8 239 2.605e-14
C276 9 239 5.64e-14
C271 14 239 5.812e-14
C270 15 239 1.2452e-13
C269 16 239 1.1722e-13
C268 17 239 1.8635e-14
C266 19 239 1.8635e-14
C265 20 239 5.529e-14
C263 22 239 2.639e-14
C261 24 239 1.4489e-13
C260 25 239 1.8635e-14
C259 26 239 4.783e-14
C258 27 239 7.476e-14
C255 30 239 6.082e-14
C254 31 239 4.595e-14
C247 38 239 7.768e-14
C243 42 239 6.876e-14
C240 45 239 6.052e-14
C237 48 239 5.482e-14
C235 50 239 7.325e-14
C234 51 239 6.05e-15
C231 53 239 9.7e-15
C228 56 239 2.1714e-13
C225 59 239 6.316e-14
C224 60 239 5.37e-14
C223 61 239 1.0516e-13
C222 62 239 8.419e-14
C221 63 239 1.8635e-14
C220 64 239 1.1774e-13
C215 69 239 1.767e-14
C213 71 239 2.596e-14
C212 72 239 2.16e-14
C211 73 239 1.0534e-13
C209 74 239 2.931e-14
C208 75 239 8.248e-14
C205 78 239 5.242e-14
C204 79 239 5.991e-14
C200 83 239 6.022e-14
C199 84 239 2.596e-14
C198 85 239 8.115e-14
C197 86 239 1.6456e-13
C196 87 239 6.21e-14
C195 88 239 2.16e-14
C194 89 239 7.76e-15
C193 90 239 2.605e-14
C192 91 239 1.3797e-13
C190 93 239 4.839e-14
C189 94 239 1.1068e-13
C188 95 239 7.666e-14
C185 98 239 5.746e-14
C181 102 239 8.08e-14
C180 103 239 1.0726e-13
C174 109 239 9.022e-14
C170 113 239 8.466e-14
C157 125 239 4.987e-14
C156 126 239 5.312e-14
C155 127 239 4.11e-15
C151 131 239 2.605e-14
C150 132 239 7.741e-14
C149 133 239 4.11e-15
C148 134 239 4.515e-14
C147 135 239 7.452e-14
C145 137 239 6.306e-14
C142 140 239 2.0905e-13
C141 141 239 5.064e-14
C137 145 239 2.2285e-13
C136 146 239 2.306e-14
C135 147 239 1.0545e-13
C134 148 239 9.058e-14
C133 149 239 8.817e-14
C130 152 239 1.1276e-13
C127 155 239 1.035e-13
C122 159 239 3.101e-13
C121 160 239 2.596e-14
C120 161 239 2.16e-14
C119 162 239 3.889e-14
C118 163 239 9.7e-15
C117 164 239 2.596e-14
C116 165 239 9.7e-15
C115 166 239 4.369e-14
C114 167 239 2.16e-14
C113 168 239 9.295e-14
C112 169 239 1.5137e-13
C110 171 239 2.596e-14
C109 172 239 2.16e-14
C108 173 239 9.7e-15
C107 174 239 1.568e-14
C106 175 239 7.689e-14
C105 176 239 5.169e-14
C104 177 239 5.965e-14
C103 178 239 2.445e-14
C102 179 239 7.43e-15
C101 180 239 1.8635e-14
C100 181 239 8.852e-14
C99 182 239 1.3034e-13
C98 183 239 2.596e-14
C97 184 239 2.16e-14
C96 185 239 7.405e-14
C95 186 239 9.7e-15
C94 187 239 2.5762e-13
C93 188 239 1.8635e-14
C92 189 239 8.7e-14
C91 190 239 6.05e-15
C86 195 239 6.05e-15
C81 199 239 5.981e-14
C78 202 239 2.605e-14
C77 203 239 1.2366e-13
C76 204 239 1.767e-14
C71 209 239 5.747e-14
C70 210 239 2.455e-14
C69 211 239 1.8454e-13
C68 212 239 4.11e-15
C67 213 239 4.123e-14
C66 214 239 1.568e-14
C63 217 239 1.0572e-13
C62 218 239 1.242e-13
C61 219 239 1.8635e-14
C60 220 239 2.4222e-13
C58 222 239 1.8635e-14
C55 225 239 1.3861e-13
C54 226 239 1.8635e-14
C52 228 239 1.3011e-13
C51 229 239 1.8635e-14
C48 232 239 9.776e-14
C47 233 239 1.568e-14
C46 234 239 5.053e-14
C45 235 239 1.8635e-14
C43 237 239 1.3313e-13
C41 239 239 3.22324e-12
C40 240 239 7.497e-14
C39 241 239 2.445e-14
C38 242 239 7.43e-15
C37 243 239 2.596e-14
C36 244 239 5.365e-14
C35 245 239 9.7e-15
C34 246 239 2.3489e-13
C33 247 239 2.16e-14
C32 248 239 7.75e-14
C31 249 239 1.6918e-13
C30 250 239 2.596e-14
C29 251 239 6.685e-14
C28 252 239 9.7e-15
C27 253 239 2.16e-14
C26 254 239 1.0338e-13
C25 255 239 1.568e-14
C24 256 239 2.8904e-13
C23 257 239 5.169e-14
C22 258 239 2.371e-13
C21 259 239 2.422e-13
C20 260 239 1.1122e-13
C19 261 239 1.1278e-13
C18 262 239 9.754e-14
C17 263 239 1.8635e-14
C15 265 239 8.413e-14
C14 266 239 2.6041e-13
C13 267 239 2.3605e-13
C12 268 239 1.0849e-13
C11 269 239 9.7e-15
C10 270 239 2.596e-14
C9 271 239 2.1135e-13
C8 272 239 2.16e-14
C7 273 239 1.4797e-13
C6 274 239 1.4742e-13
C5 275 239 2.596e-14
C4 276 239 2.16e-14
C3 277 239 5.991e-14
C2 278 239 3.33076e-12
C1 279 239 9.7e-15
.ends sum5b_cougar

