* Spice description of mul3b_cougar
* Spice driver version -1208766812
* Date ( dd/mm/yyyy hh:mm:ss ):  4/11/2020 at 11:12:56

* INTERF vdd vss x[0] x[1] x[2] y[0] y[1] y[2] z[0] z[1] z[2] z[3] z[4] z[5] 


.subckt mul3b_cougar vdd vss x[0] x[1] x[2] y[0] y[1] y[2] z[0] z[1] z[2] z[3] z[4] z[5] 
Mtr_00408 sig7 rtl_map_5 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00407 vdd u0.x1 sig1 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00406 u0.y0.xr2_x1_sig sig7 sig5 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00405 sig5 u0.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00404 sig5 sig1 u0.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00403 vdd rtl_map_5 sig5 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00402 sig16 rtl_map_4 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00401 vdd u0.y0.xr2_x1_sig sig13 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00400 sx[0] sig16 sig14 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00399 sig14 u0.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00398 sig14 sig13 sx[0] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00397 vdd rtl_map_4 sig14 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00396 z[0] sig23 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00395 vdd sx[0] sig23 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00394 cx[0] sig10 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00393 sig8 u0.x1 sig9 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00392 sig8 rtl_map_5 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00391 vdd u0.x1 sig8 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00390 sig9 rtl_map_5 sig10 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00389 sig10 rtl_map_4 sig8 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00388 sig22 rtl_map_1 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00387 vdd u3.y0.xr2_x1_sig sig20 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00386 sx[3] sig22 sig18 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00385 sig18 u3.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00384 sig18 sig20 sx[3] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00383 vdd rtl_map_1 sig18 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00382 u3.x1 sig42 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00381 vdd y[1] sig42 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 sig42 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00379 u0.x1 sig31 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00378 vdd y[0] sig31 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00377 sig31 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00376 cx[3] sig49 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00375 sig61 u3.x1 sig62 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00374 sig61 sx[1] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00373 vdd u3.x1 sig61 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00372 sig62 sx[1] sig49 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00371 sig49 rtl_map_1 sig61 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00370 sig40 cx[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00369 vdd u1.y0.xr2_x1_sig sig34 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00368 sx[1] sig40 sig60 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00367 sig60 u1.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00366 sig60 sig34 sx[1] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00365 vdd cx[0] sig60 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00364 z[1] sig58 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00363 vdd sx[3] sig58 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00362 sig57 sx[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00361 vdd u3.x1 sig55 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00360 u3.y0.xr2_x1_sig sig57 sig63 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00359 sig63 u3.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00358 sig63 sig55 u3.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00357 vdd sx[1] sig63 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00356 u1.x1 sig64 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00355 vdd y[0] sig64 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00354 sig64 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00353 u4.x1 sig74 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00352 vdd y[1] sig74 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00351 sig74 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00350 u6.x1 sig77 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00349 vdd y[2] sig77 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00348 sig77 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00347 sig84 cx[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00346 vdd u4.y0.xr2_x1_sig sig79 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00345 sx[4] sig84 sig82 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00344 sig82 u4.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00343 sig82 sig79 sx[4] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00342 vdd cx[3] sig82 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00341 cx[1] sig73 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00340 sig71 u1.x1 sig72 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00339 sig71 rtl_map_3 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00338 vdd u1.x1 sig71 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00337 sig72 rtl_map_3 sig73 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00336 sig73 cx[0] sig71 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00335 sig70 rtl_map_3 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 vdd u1.x1 sig69 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00333 u1.y0.xr2_x1_sig sig70 sig68 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00332 sig68 u1.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00331 sig68 sig69 u1.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00330 vdd rtl_map_3 sig68 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00329 sig88 sx[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00328 vdd u6.x1 sig86 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00327 u6.y0.xr2_x1_sig sig88 sig85 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00326 sig85 u6.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00325 sig85 sig86 u6.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00324 vdd sx[4] sig85 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00323 sig90 rtl_map_0 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00322 vdd u6.y0.xr2_x1_sig sig89 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00321 sx[6] sig90 sig92 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00320 sig92 u6.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00319 sig92 sig89 sx[6] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00318 vdd rtl_map_0 sig92 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00317 z[2] sig94 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00316 vdd sx[6] sig94 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00315 sig106 rtl_map_2 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00314 vdd u2.x1 sig105 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00313 u2.y0.xr2_x1_sig sig106 sig136 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00312 sig136 u2.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00311 sig136 sig105 u2.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00310 vdd rtl_map_2 sig136 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00309 cx[2] sig99 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00308 sig132 u2.x1 sig134 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00307 sig132 rtl_map_2 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00306 vdd u2.x1 sig132 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00305 sig134 rtl_map_2 sig99 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00304 sig99 cx[1] sig132 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00303 cx[4] sig118 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00302 sig141 u4.x1 sig140 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00301 sig141 sx[2] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00300 vdd u4.x1 sig141 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00299 sig140 sx[2] sig118 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00298 sig118 cx[3] sig141 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00297 sig123 sx[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00296 vdd u4.x1 sig122 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 u4.y0.xr2_x1_sig sig123 sig143 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00294 sig143 u4.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00293 sig143 sig122 u4.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00292 vdd sx[2] sig143 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00291 sig113 cx[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 vdd u2.y0.xr2_x1_sig sig114 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 sx[2] sig113 sig137 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00288 sig137 u2.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00287 sig137 sig114 sx[2] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00286 vdd cx[1] sig137 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00285 z[3] sig129 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00284 vdd sx[7] sig129 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00283 cx[6] sig127 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00282 sig147 u6.x1 sig146 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00281 sig147 sx[4] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00280 vdd u6.x1 sig147 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00279 sig146 sx[4] sig127 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00278 sig127 rtl_map_0 sig147 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00277 sig156 cx[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 vdd u5.y0.xr2_x1_sig sig152 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 sx[5] sig156 sig154 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00274 sig154 u5.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00273 sig154 sig152 sx[5] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00272 vdd cx[4] sig154 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00271 u7.x1 sig162 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00270 vdd y[2] sig162 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00269 sig162 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 u2.x1 sig150 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00267 vdd y[0] sig150 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00266 sig150 x[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00265 sig161 sx[5] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00264 vdd u7.x1 sig157 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00263 u7.y0.xr2_x1_sig sig161 sig159 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00262 sig159 u7.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00261 sig159 sig157 u7.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00260 vdd sx[5] sig159 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00259 cx[7] sig165 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00258 sig163 u7.x1 sig164 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00257 sig163 sx[5] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00256 vdd u7.x1 sig163 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00255 sig164 sx[5] sig165 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00254 sig165 cx[6] sig163 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00253 z[4] sig175 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00252 vdd sx[8] sig175 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00251 sig169 cx[6] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00250 vdd u7.y0.xr2_x1_sig sig166 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00249 sx[7] sig169 sig168 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00248 sig168 u7.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00247 sig168 sig166 sx[7] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00246 vdd cx[6] sig168 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00245 sig174 cx[7] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 vdd u8.y0.xr2_x1_sig sig170 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 sx[8] sig174 sig173 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00242 sig173 u8.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00241 sig173 sig170 sx[8] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00240 vdd cx[7] sig173 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00239 sig179 cx[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00238 vdd u5.x1 sig181 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 u5.y0.xr2_x1_sig sig179 sig202 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00236 sig202 u5.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00235 sig202 sig181 u5.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00234 vdd cx[2] sig202 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00233 u5.x1 sig187 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00232 vdd y[1] sig187 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 sig187 x[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 cx[5] sig205 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00229 sig207 u5.x1 sig208 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00228 sig207 cx[2] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00227 vdd u5.x1 sig207 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00226 sig208 cx[2] sig205 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00225 sig205 cx[4] sig207 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00224 u8.x1 sig189 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00223 vdd y[2] sig189 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00222 sig189 x[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00221 sig195 cx[5] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 vdd u8.x1 sig193 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 u8.y0.xr2_x1_sig sig195 sig213 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00218 sig213 u8.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00217 sig213 sig193 u8.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00216 vdd cx[5] sig213 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00215 z[5] sig199 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00214 vdd cx[8] sig199 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00213 cx[8] sig214 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00212 sig217 u8.x1 sig218 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00211 sig217 cx[5] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00210 vdd u8.x1 sig217 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00209 sig218 cx[5] sig214 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00208 sig214 cx[7] sig217 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00207 sig1 u0.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00206 vss rtl_map_5 sig7 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00205 sig29 sig7 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 u0.y0.xr2_x1_sig sig1 sig29 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00203 sig30 rtl_map_5 u0.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00202 vss u0.x1 sig30 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 sig13 u0.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00200 vss rtl_map_4 sig16 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00199 sig47 sig16 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 sx[0] sig13 sig47 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 sig46 rtl_map_4 sx[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 vss u0.y0.xr2_x1_sig sig46 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00195 vss sig23 z[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00194 sig23 sx[0] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00193 vss sig10 cx[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 vss rtl_map_5 sig37 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00191 sig37 u0.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00190 sig10 rtl_map_5 sig38 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00189 sig38 u0.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00188 sig37 rtl_map_4 sig10 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00187 vss vdd rtl_map_4 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00186 vss vdd rtl_map_1 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00185 vss vdd rtl_map_5 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00184 sig20 u3.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00183 vss rtl_map_1 sig22 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00182 sig53 sig22 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00181 sx[3] sig20 sig53 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 sig52 rtl_map_1 sx[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 vss u3.y0.xr2_x1_sig sig52 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00178 vss vdd rtl_map_2 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00177 sig42 x[0] sig43 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 vss sig42 u3.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 sig43 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 sig31 x[0] sig32 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 vss sig31 u0.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00172 sig32 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 vss sig49 cx[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 vss sx[1] sig48 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00169 sig48 u3.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00168 sig49 sx[1] sig50 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00167 sig50 u3.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00166 sig48 rtl_map_1 sig49 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00165 sig34 u1.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00164 vss cx[0] sig40 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00163 sig39 sig40 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 sx[1] sig34 sig39 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 sig35 cx[0] sx[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00160 vss u1.y0.xr2_x1_sig sig35 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 vss sig58 z[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 sig58 sx[3] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00157 sig55 u3.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00156 vss sx[1] sig57 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00155 sig54 sig57 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 u3.y0.xr2_x1_sig sig55 sig54 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00153 sig56 sx[1] u3.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 vss u3.x1 sig56 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 sig64 x[1] sig96 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 vss sig64 u1.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 sig96 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00148 sig74 x[1] sig109 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 vss sig74 u4.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 sig109 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00145 sig77 x[0] sig115 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00144 vss sig77 u6.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00143 sig115 y[2] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 vss vdd rtl_map_3 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00141 sig79 u4.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00140 vss cx[3] sig84 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00139 sig116 sig84 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 sx[4] sig79 sig116 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 sig117 cx[3] sx[4] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 vss u4.y0.xr2_x1_sig sig117 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 vss sig73 cx[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 vss rtl_map_3 sig108 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00133 sig108 u1.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00132 sig73 rtl_map_3 sig101 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00131 sig101 u1.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00130 sig108 cx[0] sig73 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00129 sig69 u1.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00128 vss rtl_map_3 sig70 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00127 sig100 sig70 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 u1.y0.xr2_x1_sig sig69 sig100 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 sig98 rtl_map_3 u1.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 vss u1.x1 sig98 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00123 sig86 u6.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00122 vss sx[4] sig88 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00121 sig124 sig88 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 u6.y0.xr2_x1_sig sig86 sig124 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 sig119 sx[4] u6.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 vss u6.x1 sig119 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 sig89 u6.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00116 vss rtl_map_0 sig90 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00115 sig125 sig90 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 sx[6] sig89 sig125 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 sig126 rtl_map_0 sx[6] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 vss u6.y0.xr2_x1_sig sig126 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 vss sig94 z[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 sig94 sx[6] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00109 sig105 u2.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00108 vss rtl_map_2 sig106 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 sig102 sig106 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 u2.y0.xr2_x1_sig sig105 sig102 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 sig103 rtl_map_2 u2.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 vss u2.x1 sig103 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 vss sig99 cx[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 vss rtl_map_2 sig130 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00101 sig130 u2.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00100 sig99 rtl_map_2 sig131 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00099 sig131 u2.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00098 sig130 cx[1] sig99 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00097 vss sig118 cx[4] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 vss sx[2] sig138 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00095 sig138 u4.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00094 sig118 sx[2] sig139 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00093 sig139 u4.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00092 sig138 cx[3] sig118 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00091 sig122 u4.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00090 vss sx[2] sig123 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00089 sig120 sig123 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 u4.y0.xr2_x1_sig sig122 sig120 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 sig121 sx[2] u4.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 vss u4.x1 sig121 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 sig114 u2.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00084 vss cx[1] sig113 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00083 sig110 sig113 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 sx[2] sig114 sig110 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 sig111 cx[1] sx[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 vss u2.y0.xr2_x1_sig sig111 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 vss sig129 z[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 sig129 sx[7] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00077 vss sig127 cx[6] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 vss sx[4] sig144 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00075 sig144 u6.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00074 sig127 sx[4] sig145 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00073 sig145 u6.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00072 sig144 rtl_map_0 sig127 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00071 vss vdd rtl_map_0 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00070 sig152 u5.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 vss cx[4] sig156 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00068 sig182 sig156 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 sx[5] sig152 sig182 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 sig183 cx[4] sx[5] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 vss u5.y0.xr2_x1_sig sig183 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 sig162 x[1] sig186 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 vss sig162 u7.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 sig186 y[2] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 sig150 x[2] sig177 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 vss sig150 u2.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 sig177 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 sig157 u7.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00057 vss sx[5] sig161 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 sig185 sig161 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 u7.y0.xr2_x1_sig sig157 sig185 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 sig184 sx[5] u7.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 vss u7.x1 sig184 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 vss sig165 cx[7] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 vss sx[5] sig190 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00050 sig190 u7.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00049 sig165 sx[5] sig188 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00048 sig188 u7.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00047 sig190 cx[6] sig165 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00046 vss sig175 z[4] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 sig175 sx[8] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00044 sig166 u7.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00043 vss cx[6] sig169 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00042 sig196 sig169 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 sx[7] sig166 sig196 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 sig194 cx[6] sx[7] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 vss u7.y0.xr2_x1_sig sig194 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 sig170 u8.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00037 vss cx[7] sig174 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00036 sig198 sig174 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 sx[8] sig170 sig198 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 sig197 cx[7] sx[8] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 vss u8.y0.xr2_x1_sig sig197 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 sig181 u5.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00031 vss cx[2] sig179 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00030 sig200 sig179 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 u5.y0.xr2_x1_sig sig181 sig200 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 sig201 cx[2] u5.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 vss u5.x1 sig201 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 sig187 x[2] sig209 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 vss sig187 u5.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 sig209 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 vss sig205 cx[5] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 vss cx[2] sig204 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00021 sig204 u5.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00020 sig205 cx[2] sig206 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00019 sig206 u5.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00018 sig204 cx[4] sig205 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00017 sig189 x[2] sig210 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 vss sig189 u8.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 sig210 y[2] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 sig193 u8.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 vss cx[5] sig195 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 sig211 sig195 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 u8.y0.xr2_x1_sig sig193 sig211 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 sig212 cx[5] u8.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 vss u8.x1 sig212 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 vss sig199 z[5] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 sig199 cx[8] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00006 vss sig214 cx[8] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 vss cx[5] sig215 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00004 sig215 u8.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00003 sig214 cx[5] sig216 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00002 sig216 u8.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00001 sig215 cx[7] sig214 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
C220 z[5] vss 2.659e-14
C219 cx[8] vss 5.333e-14
C217 sig217 vss 8.58e-15
C215 sig215 vss 4.11e-15
C214 sig214 vss 2.299e-14
C213 sig213 vss 9.7e-15
C207 sig207 vss 8.58e-15
C205 sig205 vss 2.299e-14
C204 sig204 vss 4.11e-15
C202 sig202 vss 9.7e-15
C199 sig199 vss 1.568e-14
C195 sig195 vss 2.596e-14
C193 sig193 vss 2.16e-14
C192 cx[5] vss 1.3096e-13
C191 u8.x1 vss 1.1131e-13
C190 sig190 vss 4.11e-15
C189 sig189 vss 1.8635e-14
C187 sig187 vss 1.8635e-14
C181 sig181 vss 2.16e-14
C180 u5.x1 vss 1.1291e-13
C179 sig179 vss 2.596e-14
C176 z[4] vss 2.371e-14
C175 sig175 vss 1.568e-14
C174 sig174 vss 2.596e-14
C173 sig173 vss 9.7e-15
C172 sx[8] vss 5.619e-14
C171 u8.y0.xr2_x1_sig vss 7.551e-14
C170 sig170 vss 2.16e-14
C169 sig169 vss 2.596e-14
C168 sig168 vss 9.7e-15
C167 cx[7] vss 1.1053e-13
C166 sig166 vss 2.16e-14
C165 sig165 vss 2.299e-14
C163 sig163 vss 8.58e-15
C162 sig162 vss 1.8635e-14
C161 sig161 vss 2.596e-14
C160 u7.x1 vss 1.1371e-13
C159 sig159 vss 9.7e-15
C158 u7.y0.xr2_x1_sig vss 8.151e-14
C157 sig157 vss 2.16e-14
C156 sig156 vss 2.596e-14
C155 u5.y0.xr2_x1_sig vss 6.231e-14
C154 sig154 vss 9.7e-15
C153 sx[5] vss 1.2222e-13
C152 sig152 vss 2.16e-14
C151 x[2] vss 1.006e-13
C150 sig150 vss 1.8635e-14
C149 sx[7] vss 7.539e-14
C148 cx[6] vss 1.0909e-13
C147 sig147 vss 8.58e-15
C144 sig144 vss 4.11e-15
C143 sig143 vss 9.7e-15
C142 cx[4] vss 1.2949e-13
C141 sig141 vss 8.58e-15
C138 sig138 vss 4.11e-15
C137 sig137 vss 9.7e-15
C136 sig136 vss 9.7e-15
C135 cx[2] vss 1.2056e-13
C132 sig132 vss 8.58e-15
C130 sig130 vss 4.11e-15
C129 sig129 vss 1.568e-14
C128 z[3] vss 2.371e-14
C127 sig127 vss 2.299e-14
C123 sig123 vss 2.596e-14
C122 sig122 vss 2.16e-14
C118 sig118 vss 2.299e-14
C114 sig114 vss 2.16e-14
C113 sig113 vss 2.596e-14
C112 sx[2] vss 1.1718e-13
C108 sig108 vss 4.11e-15
C107 u2.x1 vss 1.0883e-13
C106 sig106 vss 2.596e-14
C105 sig105 vss 2.16e-14
C104 u2.y0.xr2_x1_sig vss 5.991e-14
C99 sig99 vss 2.299e-14
C95 z[2] vss 2.371e-14
C94 sig94 vss 1.568e-14
C93 rtl_map_0 vss 9.109e-14
C92 sig92 vss 9.7e-15
C91 sx[6] vss 5.619e-14
C90 sig90 vss 2.596e-14
C89 sig89 vss 2.16e-14
C88 sig88 vss 2.596e-14
C87 u6.y0.xr2_x1_sig vss 5.751e-14
C86 sig86 vss 2.16e-14
C85 sig85 vss 9.7e-15
C84 sig84 vss 2.596e-14
C83 u4.y0.xr2_x1_sig vss 6.351e-14
C82 sig82 vss 9.7e-15
C81 sx[4] vss 1.1798e-13
C80 y[2] vss 1.5555e-13
C79 sig79 vss 2.16e-14
C78 u6.x1 vss 1.2467e-13
C77 sig77 vss 1.8635e-14
C76 cx[1] vss 1.2021e-13
C75 u4.x1 vss 1.1131e-13
C74 sig74 vss 1.8635e-14
C73 sig73 vss 2.299e-14
C71 sig71 vss 8.58e-15
C70 sig70 vss 2.596e-14
C69 sig69 vss 2.16e-14
C68 sig68 vss 9.7e-15
C67 u1.x1 vss 1.1331e-13
C66 rtl_map_3 vss 1.0632e-13
C65 x[1] vss 1.1572e-13
C64 sig64 vss 1.8635e-14
C63 sig63 vss 9.7e-15
C61 sig61 vss 8.58e-15
C60 sig60 vss 9.7e-15
C59 z[1] vss 2.659e-14
C58 sig58 vss 1.568e-14
C57 sig57 vss 2.596e-14
C55 sig55 vss 2.16e-14
C51 cx[3] vss 1.0669e-13
C49 sig49 vss 2.299e-14
C48 sig48 vss 4.11e-15
C45 u3.x1 vss 1.1251e-13
C44 y[1] vss 1.5315e-13
C42 sig42 vss 1.8635e-14
C41 sx[1] vss 1.3182e-13
C40 sig40 vss 2.596e-14
C37 sig37 vss 4.11e-15
C36 u1.y0.xr2_x1_sig vss 6.591e-14
C34 sig34 vss 2.16e-14
C33 y[0] vss 1.5867e-13
C31 sig31 vss 1.8635e-14
C28 x[0] vss 1.0804e-13
C27 rtl_map_2 vss 1.2312e-13
C25 vss vss 2.4434e-12
C24 z[0] vss 2.659e-14
C23 sig23 vss 1.568e-14
C22 sig22 vss 2.596e-14
C21 u3.y0.xr2_x1_sig vss 5.751e-14
C20 sig20 vss 2.16e-14
C19 sx[3] vss 6.579e-14
C18 sig18 vss 9.7e-15
C17 rtl_map_1 vss 1.0589e-13
C16 sig16 vss 2.596e-14
C15 sx[0] vss 7.779e-14
C14 sig14 vss 9.7e-15
C13 sig13 vss 2.16e-14
C12 cx[0] vss 9.949e-14
C11 rtl_map_4 vss 9.901e-14
C10 sig10 vss 2.299e-14
C8 sig8 vss 8.58e-15
C7 sig7 vss 2.596e-14
C6 u0.y0.xr2_x1_sig vss 8.391e-14
C5 sig5 vss 9.7e-15
C4 rtl_map_5 vss 1.2112e-13
C3 u0.x1 vss 1.1491e-13
C2 vdd vss 2.56548e-12
C1 sig1 vss 2.16e-14
.ends mul3b_cougar

