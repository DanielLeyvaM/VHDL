* Spice description of mul4b_cougar
* Spice driver version -1209393500
* Date ( dd/mm/yyyy hh:mm:ss ): 28/10/2020 at 15:21:13

* INTERF vdd vss x[0] x[1] x[2] x[3] y[0] y[1] y[2] y[3] z[0] z[1] z[2] z[3] 
* INTERF z[4] z[5] z[6] z[7] 


.subckt mul4b_cougar 622 578 573 595 473 528 510 604 614 566 579 456 368 512 377 166 98 24 
* NET 10 = not_aux32
* NET 11 = na2_x1_15_sig
* NET 13 = on12_x1_sig
* NET 17 = na2_x1_14_sig
* NET 19 = na2_x1_12_sig
* NET 22 = na4_x1_sig
* NET 24 = z[7]
* NET 28 = a2_x2_8_sig
* NET 40 = mbk_buf_not_aux21
* NET 44 = na2_x1_11_sig
* NET 45 = o2_x2_sig
* NET 51 = aux39
* NET 53 = nao22_x1_7_sig
* NET 55 = na3_x1_9_sig
* NET 56 = an12_x1_sig
* NET 59 = na3_x1_8_sig
* NET 60 = na3_x1_7_sig
* NET 64 = na2_x1_10_sig
* NET 65 = nao22_x1_8_sig
* NET 67 = ao22_x2_8_sig
* NET 70 = oa2a22_x2_3_sig
* NET 71 = not_aux47
* NET 75 = aux21
* NET 77 = mbk_buf_aux21
* NET 79 = na2_x1_13_sig
* NET 80 = not_aux21
* NET 98 = z[6]
* NET 101 = oa2a2a23_x2_sig
* NET 103 = ao22_x2_6_sig
* NET 107 = aux45
* NET 108 = a3_x2_5_sig
* NET 114 = ao22_x2_7_sig
* NET 118 = a2_x2_7_sig
* NET 126 = nxr2_x1_3_sig
* NET 128 = na2_x1_9_sig
* NET 138 = aux43
* NET 141 = not_aux31
* NET 144 = na2_x1_6_sig
* NET 150 = nxr2_x1_2_sig
* NET 152 = aux0
* NET 155 = not_aux28
* NET 156 = ao22_x2_5_sig
* NET 159 = aux30
* NET 160 = noa22_x1_5_sig
* NET 164 = aux46
* NET 166 = z[5]
* NET 168 = oa2ao222_x2_3_sig
* NET 174 = no2_x1_6_sig
* NET 175 = inv_x2_7_sig
* NET 176 = aux32
* NET 180 = oa2ao222_x2_4_sig
* NET 181 = mx3_x2_3_sig
* NET 189 = nao2o22_x1_sig
* NET 192 = not_aux15
* NET 195 = a2_x2_5_sig
* NET 196 = not_aux33
* NET 219 = oa22_x2_3_sig
* NET 223 = na2_x1_8_sig
* NET 224 = aux2
* NET 225 = ao22_x2_4_sig
* NET 226 = noa22_x1_7_sig
* NET 230 = oa2ao222_x2_2_sig
* NET 231 = a2_x2_4_sig
* NET 235 = inv_x2_5_sig
* NET 236 = not_aux44
* NET 239 = mx3_x2_4_sig
* NET 244 = xr2_x1_8_sig
* NET 247 = inv_x2_6_sig
* NET 251 = not_aux20
* NET 252 = aux12
* NET 255 = aux27
* NET 261 = a3_x2_6_sig
* NET 262 = not_y[0]
* NET 265 = na3_x1_10_sig
* NET 270 = xr2_x1_sig
* NET 275 = no3_x1_sig
* NET 280 = not_aux18
* NET 286 = inv_x2_4_sig
* NET 290 = na2_x1_3_sig
* NET 293 = aux16
* NET 296 = not_aux38
* NET 299 = na2_x1_sig
* NET 308 = not_aux2
* NET 309 = aux1
* NET 315 = a3_x2_4_sig
* NET 319 = na3_x1_4_sig
* NET 320 = oa22_x2_2_sig
* NET 321 = na2_x1_4_sig
* NET 331 = xr2_x1_2_sig
* NET 334 = not_aux1
* NET 336 = noa22_x1_sig
* NET 340 = not_y[3]
* NET 341 = o3_x2_3_sig
* NET 343 = na3_x1_6_sig
* NET 344 = noa22_x1_6_sig
* NET 345 = na2_x1_7_sig
* NET 347 = aux17
* NET 349 = not_y[2]
* NET 352 = o3_x2_2_sig
* NET 353 = noa22_x1_4_sig
* NET 355 = not_aux13
* NET 361 = aux10
* NET 363 = mbk_buf_aux10
* NET 364 = na3_x1_sig
* NET 366 = not_aux22
* NET 368 = z[2]
* NET 371 = not_aux40
* NET 377 = z[4]
* NET 385 = aux41
* NET 390 = oa22_x2_sig
* NET 399 = not_aux0
* NET 402 = a2_x2_sig
* NET 407 = aux40
* NET 410 = not_aux3
* NET 411 = mbk_buf_not_aux40
* NET 412 = na3_x1_3_sig
* NET 415 = oa2a22_x2_2_sig
* NET 420 = mx3_x2_sig
* NET 421 = oa2ao222_x2_sig
* NET 431 = ao22_x2_3_sig
* NET 432 = no2_x1_2_sig
* NET 436 = a2_x2_2_sig
* NET 439 = xr2_x1_6_sig
* NET 448 = not_aux10
* NET 452 = na2_x1_2_sig
* NET 453 = mbk_buf_not_aux22
* NET 455 = noa22_x1_2_sig
* NET 456 = z[1]
* NET 458 = aux42
* NET 460 = a2_x2_3_sig
* NET 461 = not_aux42
* NET 464 = nao22_x1_5_sig
* NET 465 = no2_x1_4_sig
* NET 467 = nao22_x1_6_sig
* NET 468 = noa22_x1_3_sig
* NET 469 = a3_x2_3_sig
* NET 470 = na3_x1_5_sig
* NET 472 = not_x[3]
* NET 473 = x[2]
* NET 477 = not_aux24
* NET 478 = nao22_x1_4_sig
* NET 480 = mbk_buf_not_aux25
* NET 482 = not_aux23
* NET 483 = mx3_x2_2_sig
* NET 485 = inv_x2_2_sig
* NET 492 = not_aux25
* NET 493 = inv_x2_3_sig
* NET 510 = y[0]
* NET 512 = z[3]
* NET 520 = not_aux12
* NET 521 = no2_x1_3_sig
* NET 523 = xr2_x1_5_sig
* NET 528 = x[3]
* NET 530 = xr2_x1_3_sig
* NET 534 = oa2a22_x2_sig
* NET 541 = a3_x2_2_sig
* NET 545 = not_aux6
* NET 548 = aux11
* NET 549 = xr2_x1_4_sig
* NET 559 = xr2_x1_7_sig
* NET 564 = aux4
* NET 566 = y[3]
* NET 573 = x[0]
* NET 574 = no2_x1_sig
* NET 577 = not_x[0]
* NET 578 = vss
* NET 579 = z[0]
* NET 582 = na2_x1_5_sig
* NET 583 = not_aux5
* NET 584 = nao22_x1_sig
* NET 586 = not_x[2]
* NET 587 = inv_x2_sig
* NET 589 = a3_x2_sig
* NET 590 = aux7
* NET 592 = nao22_x1_3_sig
* NET 593 = nao22_x1_2_sig
* NET 594 = na3_x1_2_sig
* NET 595 = x[1]
* NET 599 = o3_x2_sig
* NET 600 = ao22_x2_2_sig
* NET 604 = y[1]
* NET 605 = not_aux8
* NET 606 = not_aux9
* NET 608 = ao22_x2_sig
* NET 611 = not_x[1]
* NET 612 = a2_x2_6_sig
* NET 614 = y[2]
* NET 616 = xr2_x1_9_sig
* NET 619 = nxr2_x1_sig
* NET 620 = not_y[1]
* NET 621 = not_aux4
* NET 622 = vdd
* NET 623 = no2_x1_5_sig
Mtr_01208 615 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01207 622 623 618 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01206 616 615 617 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01205 617 623 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01204 617 618 616 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01203 622 614 617 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01202 624 621 623 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01201 622 620 624 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01200 612 613 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01199 622 611 613 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01198 613 616 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01197 622 604 598 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01196 598 595 596 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01195 596 621 597 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01194 599 597 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01193 622 609 608 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01192 609 606 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01191 622 619 610 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01190 610 620 609 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01189 581 621 580 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01188 622 595 581 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01187 583 580 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01186 603 605 607 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01185 622 604 603 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01184 606 607 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01183 622 601 600 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01182 601 599 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01181 622 606 602 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01180 602 611 601 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01179 622 586 593 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01178 588 587 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01177 593 589 588 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01176 622 583 584 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01175 585 611 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01174 584 608 585 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01173 622 592 594 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01172 594 593 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01171 594 600 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01170 622 590 591 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01169 589 591 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01168 622 604 591 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01167 591 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01166 620 604 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01165 587 583 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01164 582 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01163 622 595 582 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01162 564 567 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01161 622 573 567 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01160 567 566 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01159 622 554 504 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01158 504 557 605 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01157 504 564 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01156 605 614 504 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01155 622 564 557 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01154 554 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01153 621 564 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01152 577 573 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01151 622 571 507 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01150 507 576 619 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01149 507 574 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01148 619 614 507 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01147 622 574 576 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01146 571 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01145 558 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01144 622 564 561 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01143 559 558 505 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01142 505 564 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01141 505 561 559 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01140 622 604 505 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01139 590 545 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01138 622 621 590 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01137 506 577 574 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01136 622 566 506 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01135 498 520 521 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01134 622 582 498 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01133 501 549 537 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01132 501 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01131 622 590 501 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01130 537 611 501 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01129 534 537 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01128 547 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01127 622 548 551 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01126 549 547 503 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01125 503 548 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01124 503 551 549 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01123 622 604 503 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01122 622 541 592 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01121 502 545 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01120 592 611 502 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01119 579 508 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01118 622 573 508 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01117 508 510 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01116 522 528 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01115 622 584 525 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01114 523 522 499 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01113 499 584 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01112 499 525 523 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01111 622 528 499 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01110 497 514 518 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01109 622 511 495 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01108 494 510 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01107 518 594 494 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01106 495 523 497 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01105 496 530 495 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01104 518 586 496 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01103 512 518 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01102 514 586 622 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01101 622 510 511 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01100 532 528 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01099 622 534 533 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01098 530 532 500 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01097 500 534 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01096 500 533 530 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01095 622 528 500 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01094 472 528 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01093 490 487 489 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01092 622 486 491 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01091 484 611 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01090 489 520 484 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01089 491 493 490 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01088 488 485 491 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01087 489 620 488 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01086 483 489 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01085 487 620 622 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01084 622 611 486 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01083 480 481 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01082 622 492 481 622 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01081 622 477 478 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01080 479 480 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01079 478 620 479 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01078 493 492 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01077 622 621 474 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01076 541 474 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01075 622 604 474 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01074 474 473 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01073 475 482 476 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01072 622 604 475 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01071 477 476 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01070 485 482 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01069 482 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01068 622 621 482 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01067 622 467 470 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01066 470 464 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01065 470 468 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01064 622 520 471 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01063 469 471 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01062 622 604 471 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01061 471 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01060 622 472 467 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01059 466 465 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01058 467 469 466 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01057 622 528 464 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01056 463 521 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01055 464 460 463 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01054 460 459 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01053 622 458 459 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01052 459 605 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01051 461 458 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01050 457 620 458 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01049 622 595 457 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01048 462 605 465 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01047 622 461 462 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01046 622 620 396 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01045 455 452 396 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01044 396 453 455 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01043 436 435 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01042 622 611 435 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01041 435 559 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01040 392 443 446 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01039 622 440 393 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01038 391 472 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01037 446 483 391 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01036 393 439 392 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01035 394 478 393 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01034 446 595 394 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01033 420 446 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01032 443 595 622 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01031 622 472 440 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01030 452 448 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01029 622 577 452 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01028 622 428 431 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01027 428 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01026 622 455 383 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01025 383 432 428 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01024 421 433 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01023 388 436 386 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01022 388 385 622 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01021 622 390 388 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01020 386 431 433 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01019 433 528 388 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01018 379 419 423 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01017 622 414 380 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01016 376 510 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01015 423 415 376 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01014 380 421 379 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01013 378 420 380 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01012 423 586 378 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01011 377 423 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01010 419 586 622 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01009 622 510 414 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_01008 375 470 409 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01007 375 586 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01006 622 412 375 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01005 409 473 375 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01004 415 409 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01003 381 611 385 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01002 622 528 381 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01001 382 577 548 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01000 622 448 382 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00999 411 406 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00998 622 371 406 622 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00997 372 411 432 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00996 622 410 372 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00995 370 448 407 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00994 622 604 370 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00993 371 407 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00992 397 399 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00991 622 402 398 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00990 456 397 369 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00989 369 402 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00988 369 398 456 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00987 622 399 369 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00986 402 401 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00985 622 595 401 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00984 401 510 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00983 453 367 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00982 622 366 367 622 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00981 622 361 448 622 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_00980 448 361 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00979 622 545 364 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00978 364 363 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00977 364 620 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00976 358 566 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00975 622 614 360 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00974 361 358 359 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00973 359 614 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00972 359 360 361 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00971 622 566 359 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00970 363 362 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00969 622 361 362 622 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00968 356 548 357 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00967 622 520 356 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00966 355 357 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00965 622 611 354 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00964 353 352 354 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00963 354 477 353 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00962 351 349 350 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00961 622 573 351 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00960 545 350 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00959 492 365 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00958 622 545 365 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00957 365 366 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00956 345 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00955 622 347 345 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00954 622 341 343 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00953 343 345 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00952 343 411 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00951 622 371 346 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00950 344 577 346 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00949 346 349 344 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00948 348 349 347 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00947 622 604 348 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00946 410 337 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00945 622 349 337 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00944 337 573 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00943 622 461 339 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00942 339 410 338 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00941 338 340 342 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00940 341 342 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00939 622 410 335 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00938 336 577 335 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00937 335 334 336 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00936 330 473 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00935 622 336 332 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00934 331 330 333 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00933 333 336 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00932 333 332 331 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00931 622 473 333 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00930 622 328 296 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00929 328 364 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00928 622 520 295 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00927 295 299 328 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00926 321 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00925 622 293 321 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00924 622 325 390 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00923 291 293 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00922 291 290 325 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00921 325 604 291 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00920 299 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00919 622 614 299 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00918 622 355 319 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00917 319 385 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00916 319 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00915 622 319 412 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00914 412 320 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00913 412 321 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00912 622 620 282 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00911 282 448 281 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00910 281 308 317 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00909 352 317 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00908 622 322 320 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00907 288 286 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00906 288 355 322 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00905 322 595 288 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00904 622 595 265 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00903 265 586 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00902 265 573 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00901 622 611 274 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00900 273 448 275 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00899 274 347 273 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00898 622 315 276 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00897 468 347 276 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00896 276 611 468 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00895 622 620 316 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00894 315 316 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00893 622 280 316 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00892 316 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00891 622 265 302 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00890 261 302 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00889 622 262 302 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00888 302 334 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00887 309 312 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00886 622 595 312 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00885 312 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00884 259 331 300 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00883 259 262 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00882 622 270 259 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00881 300 510 259 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00880 368 300 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00879 334 309 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00878 306 308 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00877 622 309 307 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00876 270 306 268 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00875 268 309 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00874 268 307 270 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00873 622 308 268 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00872 622 621 255 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00871 253 573 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00870 255 448 253 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00869 254 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00868 622 255 257 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00867 439 254 256 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00866 256 255 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00865 256 257 439 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00864 622 604 256 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00863 238 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00862 622 520 241 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00861 244 238 240 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00860 240 520 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00859 240 241 244 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00858 622 604 240 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00857 252 566 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00856 622 577 252 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00855 290 251 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00854 622 252 290 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00853 622 227 225 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00852 227 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00851 622 344 228 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00850 228 226 227 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00849 245 242 248 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00848 622 243 249 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00847 246 611 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00846 248 244 246 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00845 249 255 245 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00844 250 247 249 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00843 248 620 250 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00842 239 248 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00841 242 620 622 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00840 622 611 243 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00839 235 236 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00838 622 385 236 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00837 236 237 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00836 622 621 237 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00835 231 229 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00834 622 611 229 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00833 229 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00832 247 280 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00831 230 232 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00830 234 231 233 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00829 234 614 622 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00828 622 235 234 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00827 233 353 232 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00826 232 528 234 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00825 622 620 220 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00824 226 219 220 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00823 220 621 226 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00822 280 448 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00821 622 224 280 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00820 262 510 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00819 308 224 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00818 224 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00817 622 573 224 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00816 223 611 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00815 622 224 223 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00814 622 221 219 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00813 222 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00812 222 577 221 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00811 221 340 222 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00810 151 251 197 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00809 622 620 151 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00808 196 197 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00807 195 194 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00806 622 192 194 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00805 194 196 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00804 586 473 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00803 622 349 142 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00802 142 566 143 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00801 143 577 191 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00800 251 191 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00799 180 178 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00798 133 612 132 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00797 133 175 622 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00796 622 176 133 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00795 132 225 178 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00794 178 528 133 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00793 175 236 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00792 136 188 185 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00791 622 183 137 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00790 134 473 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00789 185 180 134 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00788 137 239 136 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00787 135 189 137 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00786 185 528 135 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00785 181 185 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00784 188 528 622 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00783 622 473 183 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00782 145 192 293 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00781 622 604 145 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00780 189 195 140 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00779 140 595 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00778 139 611 189 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00777 622 296 139 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00776 122 170 172 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00775 622 167 123 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00774 119 262 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00773 172 181 119 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00772 123 168 122 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00771 121 230 123 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00770 172 473 121 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00769 166 172 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00768 170 473 622 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00767 622 262 167 622 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00766 127 296 174 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00765 622 595 127 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00764 116 472 164 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00763 622 473 116 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00762 168 163 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00761 113 159 112 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00760 113 528 622 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00759 622 343 113 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00758 112 160 163 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00757 163 472 113 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00756 155 153 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00755 622 399 153 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00754 153 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00753 622 155 105 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00752 106 595 159 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00751 105 340 106 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00750 622 157 156 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00749 157 164 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00748 622 275 110 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00747 110 159 157 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00746 399 152 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00745 622 611 146 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00744 160 144 146 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00743 146 141 160 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00742 520 252 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00741 144 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00740 622 150 144 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00739 622 147 149 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00738 149 148 150 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00737 149 252 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00736 150 614 149 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00735 622 252 148 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00734 147 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00733 286 138 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00732 340 566 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00731 622 566 340 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00730 622 566 340 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00729 340 566 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00728 131 308 130 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00727 622 340 131 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00726 192 130 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00725 176 620 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00724 622 349 176 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00723 118 120 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00722 622 595 120 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00721 120 126 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00720 622 115 114 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00719 115 528 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00718 622 118 117 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00717 117 174 115 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00716 622 124 125 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00715 125 129 126 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00714 125 128 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00713 126 614 125 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00712 622 128 129 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00711 124 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00710 128 620 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00709 622 520 128 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00708 622 104 103 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00707 104 473 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00706 622 114 109 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00705 109 108 104 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00704 622 223 111 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00703 108 111 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00702 622 107 111 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00701 111 176 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00700 152 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00699 622 573 152 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00698 98 99 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00697 102 156 100 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00696 102 262 622 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00695 622 101 102 622 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00694 100 103 99 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00693 99 510 102 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00692 77 76 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00691 622 75 76 622 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00690 79 141 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00689 622 196 79 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00688 41 577 81 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00687 622 80 41 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00686 366 81 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00685 622 69 67 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00684 69 611 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00683 622 573 35 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00682 35 620 69 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00681 36 340 75 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00680 622 614 36 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00679 44 349 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00678 622 152 44 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00677 71 48 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00676 622 152 48 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00675 48 611 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00674 37 71 74 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00673 37 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00672 622 79 37 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00671 74 77 37 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00670 70 74 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00669 101 62 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00668 622 55 31 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00667 31 56 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00666 31 70 32 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00665 32 528 31 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00664 62 473 32 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00663 32 64 62 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00662 54 164 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00661 622 54 30 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00660 30 340 56 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00659 622 586 53 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00658 29 71 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00657 53 349 29 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00656 51 620 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00655 622 577 51 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00654 64 59 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00653 622 60 64 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00652 26 340 107 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00651 622 528 26 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00650 622 473 65 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00649 33 614 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00648 65 67 33 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00647 622 44 60 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00646 60 45 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00645 60 107 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00644 23 155 42 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00643 622 595 23 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00642 45 42 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00641 40 39 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00640 622 80 39 622 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00639 349 614 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00638 21 40 38 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00637 622 604 21 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00636 141 38 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00635 80 75 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00634 138 34 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00633 622 604 34 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00632 34 528 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00631 10 176 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00630 19 566 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00629 622 611 19 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00628 622 138 59 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00627 59 19 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00626 59 614 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00625 11 10 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00624 622 611 11 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00623 17 604 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00622 622 349 17 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00621 28 27 622 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00620 622 566 27 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00619 27 528 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00618 622 17 55 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00617 55 51 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00616 55 595 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00615 611 595 622 622 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00614 622 22 25 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00613 24 65 25 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00612 25 261 24 622 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00611 622 349 13 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00610 13 15 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00609 622 51 15 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00608 622 11 22 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00607 22 28 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00606 622 53 22 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00605 22 13 622 622 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00604 618 623 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00603 578 614 615 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00602 569 615 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00601 616 618 569 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00600 572 614 616 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00599 578 623 572 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00598 623 620 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00597 578 621 623 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00596 613 616 565 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00595 578 613 612 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00594 565 611 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00593 597 621 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00592 597 604 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00591 578 595 597 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00590 578 597 599 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00589 609 619 563 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00588 563 620 609 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00587 578 606 563 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00586 608 609 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00585 583 580 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00584 580 595 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00583 578 621 580 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00582 606 607 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00581 607 604 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00580 578 605 607 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00579 601 606 555 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00578 555 611 601 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00577 578 599 555 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00576 600 601 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00575 535 587 593 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00574 593 589 535 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00573 535 586 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00572 527 611 584 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00571 584 608 527 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00570 527 583 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00569 578 600 544 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00568 544 592 542 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00567 542 593 594 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00566 578 591 589 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00565 539 590 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00564 540 595 539 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00563 591 604 540 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00562 578 604 620 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00561 578 583 587 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00560 578 604 519 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00559 519 595 582 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00558 567 566 568 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00557 578 567 564 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00556 568 573 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00555 578 564 556 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00554 556 554 605 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00553 605 557 553 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00552 553 614 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00551 578 614 554 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00550 557 564 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00549 578 564 621 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00548 578 573 577 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00547 578 574 575 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00546 575 571 619 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00545 619 576 570 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00544 570 614 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00543 578 614 571 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00542 576 574 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00541 561 564 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00540 578 604 558 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00539 562 558 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00538 559 561 562 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00537 560 604 559 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00536 578 564 560 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00535 578 545 543 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00534 543 621 590 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00533 574 566 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00532 578 577 574 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00531 521 582 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00530 578 520 521 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00529 538 549 537 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00528 578 611 538 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00527 536 595 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00526 537 590 536 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00525 578 537 534 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00524 551 548 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00523 578 604 547 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00522 552 547 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00521 549 551 552 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00520 550 604 549 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00519 578 548 550 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00518 546 545 592 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00517 592 611 546 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00516 546 541 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00515 508 510 509 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00514 578 508 579 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00513 509 573 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00512 525 584 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00511 578 528 522 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00510 526 522 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00509 523 525 526 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00508 524 528 523 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00507 578 584 524 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00506 578 586 514 578 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00505 511 510 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00504 516 523 515 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00503 515 586 518 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00502 518 514 517 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00501 517 530 516 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00500 578 510 516 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00499 513 511 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00498 518 594 513 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00497 578 518 512 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00496 533 534 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00495 578 528 532 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00494 529 532 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00493 530 533 529 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00492 531 528 530 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00491 578 534 531 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00490 578 528 472 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00489 578 620 487 578 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00488 486 611 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00487 449 493 450 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00486 450 620 489 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00485 489 487 451 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00484 451 485 449 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00483 578 611 449 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00482 447 486 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00481 489 520 447 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00480 578 489 483 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00479 578 481 480 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00478 481 492 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00477 438 480 478 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00476 478 620 438 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00475 438 477 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00474 578 492 493 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00473 578 474 541 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00472 429 621 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00471 430 473 429 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00470 474 604 430 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00469 477 476 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00468 476 604 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00467 578 482 476 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00466 578 482 485 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00465 578 614 434 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00464 434 621 482 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00463 578 468 418 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00462 418 467 417 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00461 417 464 470 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00460 578 471 469 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00459 426 520 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00458 427 595 426 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00457 471 604 427 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00456 413 465 467 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00455 467 469 413 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00454 413 472 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00453 408 521 464 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00452 464 460 408 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00451 408 528 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00450 459 605 404 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00449 578 459 460 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00448 404 458 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00447 578 458 461 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00446 458 595 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00445 578 620 458 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00444 465 461 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00443 578 605 465 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00442 578 452 454 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00441 454 453 455 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00440 455 620 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00439 435 559 437 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00438 578 435 436 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00437 437 611 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00436 578 595 443 578 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00435 440 472 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00434 444 439 442 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00433 442 595 446 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00432 446 443 445 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00431 445 478 444 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00430 578 472 444 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00429 441 440 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00428 446 483 441 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00427 578 446 420 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00426 578 448 395 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00425 395 577 452 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00424 428 455 384 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00423 384 432 428 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00422 578 595 384 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00421 431 428 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00420 578 433 421 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00419 578 431 387 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00418 387 436 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00417 433 385 389 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00416 389 390 578 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00415 387 528 433 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00414 578 586 419 578 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00413 414 510 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00412 424 421 422 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00411 422 586 423 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00410 423 419 425 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00409 425 420 424 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00408 578 510 424 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00407 416 414 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00406 423 415 416 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00405 578 423 377 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00404 373 470 409 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00403 578 473 373 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00402 374 586 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00401 409 412 374 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00400 578 409 415 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00399 385 528 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00398 578 611 385 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00397 548 448 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00396 578 577 548 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00395 578 406 411 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00394 406 371 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00393 432 410 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00392 578 411 432 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00391 407 604 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00390 578 448 407 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00389 578 407 371 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00388 398 402 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00387 578 399 397 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00386 400 397 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00385 456 398 400 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 403 399 456 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00383 578 402 403 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 401 510 405 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 578 401 402 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 405 595 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00379 578 367 453 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00378 367 366 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00377 578 361 448 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00376 448 361 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00375 578 620 327 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00374 327 545 326 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00373 326 363 364 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00372 360 614 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00371 578 566 358 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00370 324 358 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00369 361 360 324 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00368 323 566 361 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00367 578 614 323 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00366 578 362 363 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00365 362 361 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00364 355 357 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00363 357 520 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00362 578 548 357 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00361 578 352 318 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00360 318 477 353 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00359 353 611 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00358 545 350 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00357 350 573 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00356 578 349 350 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00355 365 366 329 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00354 578 365 492 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00353 329 545 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00352 578 595 314 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00351 314 347 345 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00350 578 411 311 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00349 311 341 310 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00348 310 345 343 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00347 578 577 313 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00346 313 349 344 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00345 344 371 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00344 347 604 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00343 578 349 347 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00342 337 573 305 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00341 578 337 410 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00340 305 349 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00339 342 340 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00338 342 461 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00337 578 410 342 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00336 578 342 341 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00335 578 577 304 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 304 334 336 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00333 336 410 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00332 332 336 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00331 578 473 330 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00330 301 330 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00329 331 332 301 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00328 303 473 331 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00327 578 336 303 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00326 328 520 297 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00325 297 299 328 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00324 578 364 297 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00323 296 328 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00322 578 595 294 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00321 294 293 321 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00320 390 325 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00319 578 293 325 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00318 292 290 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00317 325 604 292 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00316 578 604 298 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00315 298 614 299 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00314 578 604 284 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00313 284 355 283 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00312 283 385 319 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00311 578 321 287 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00310 287 319 285 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00309 285 320 412 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00308 317 308 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00307 317 620 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00306 578 448 317 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00305 578 317 352 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00304 320 322 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 578 286 322 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00302 289 355 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00301 322 595 289 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00300 578 573 266 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00299 266 595 267 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00298 267 586 265 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00297 578 347 275 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00296 275 611 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00295 275 448 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00294 578 347 277 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 277 611 468 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 468 315 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 578 316 315 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 279 620 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 278 595 279 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00288 316 280 278 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00287 578 302 261 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00286 263 265 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00285 264 334 263 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00284 302 262 264 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00283 312 604 272 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00282 578 312 309 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 272 595 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 260 331 300 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00279 578 510 260 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00278 258 262 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00277 300 270 258 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00276 578 300 368 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 578 309 334 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 307 309 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00273 578 308 306 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00272 269 306 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00271 270 307 269 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00270 271 308 270 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00269 578 309 271 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 216 573 255 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 255 448 216 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00266 216 621 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00265 257 255 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00264 578 604 254 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00263 218 254 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 439 257 218 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 217 604 439 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 578 255 217 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00259 241 520 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00258 578 604 238 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00257 208 238 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00256 244 241 208 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00255 209 604 244 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00254 578 520 209 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00253 578 566 214 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00252 214 577 252 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00251 578 251 215 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00250 215 252 290 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00249 227 344 203 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00248 203 226 227 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00247 578 595 203 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00246 225 227 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00245 578 620 242 578 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00244 243 611 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00243 212 255 211 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00242 211 620 248 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00241 248 242 213 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00240 213 247 212 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00239 578 611 212 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00238 210 243 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00237 248 244 210 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00236 578 248 239 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00235 578 236 235 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 237 621 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00233 207 385 236 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 578 237 207 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 229 614 204 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 578 229 231 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 204 611 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00228 578 280 247 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00227 578 232 230 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00226 578 353 206 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00225 206 231 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00224 232 614 205 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00223 205 235 578 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00222 206 528 232 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00221 578 219 198 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 198 621 226 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 226 620 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 578 448 202 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 202 224 280 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 578 510 262 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00215 578 224 308 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00214 578 614 200 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 200 573 224 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 578 611 201 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 201 224 223 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00210 219 221 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00209 578 614 221 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00208 199 577 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00207 221 340 199 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00206 196 197 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00205 197 620 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00204 578 251 197 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00203 194 196 193 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00202 578 194 195 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 193 192 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 578 473 586 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 191 577 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00198 191 349 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00197 578 566 191 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00196 578 191 251 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00195 578 178 180 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00194 578 225 179 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00193 179 612 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00192 178 175 177 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00191 177 176 578 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00190 179 528 178 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00189 578 236 175 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00188 578 528 188 578 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00187 183 473 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00186 186 239 184 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00185 184 528 185 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00184 185 188 187 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00183 187 189 186 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00182 578 473 186 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00181 182 183 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00180 185 180 182 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00179 578 185 181 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00178 293 604 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00177 578 192 293 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00176 578 296 190 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 190 611 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 189 195 190 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 190 595 189 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00172 578 473 170 578 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00171 167 262 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00170 171 168 173 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00169 173 473 172 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00168 172 170 169 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00167 169 230 171 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00166 578 262 171 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00165 165 167 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00164 172 181 165 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00163 578 172 166 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 174 595 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00161 578 296 174 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00160 164 473 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00159 578 472 164 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00158 578 163 168 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00157 578 160 161 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00156 161 159 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00155 163 528 162 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00154 162 343 578 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00153 161 472 163 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00152 153 614 154 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 578 153 155 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 154 399 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 578 340 159 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00148 159 155 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00147 159 595 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00146 157 275 158 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00145 158 159 157 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00144 578 164 158 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00143 156 157 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 578 152 399 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 578 144 95 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 95 141 160 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 160 611 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 578 252 520 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 578 604 94 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 94 150 144 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 578 252 97 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 97 147 150 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00133 150 148 96 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00132 96 614 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00131 578 614 147 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00130 148 252 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00129 578 138 286 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 578 566 340 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00127 340 566 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 578 566 340 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 340 566 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 192 130 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00123 130 340 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00122 578 308 130 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00121 578 620 88 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 88 349 176 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 120 126 90 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 578 120 118 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 90 595 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 115 118 89 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00115 89 174 115 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00114 578 528 89 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00113 114 115 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 578 128 92 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 92 124 126 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 126 129 91 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 91 614 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 578 614 124 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 129 128 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00106 578 620 93 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 93 520 128 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 104 114 87 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00103 87 108 104 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00102 578 473 87 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00101 103 104 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 578 111 108 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 85 223 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00098 86 176 85 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 111 107 86 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 578 604 82 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 82 573 152 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 578 99 98 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 578 103 83 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00092 83 156 578 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00091 99 262 84 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00090 84 101 578 578 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00089 83 510 99 578 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00088 578 76 77 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 76 75 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00086 578 141 78 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 78 196 79 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00084 366 81 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 81 80 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00082 578 577 81 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00081 69 573 68 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00080 68 620 69 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00079 578 611 68 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00078 67 69 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 75 614 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00076 578 340 75 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00075 578 349 43 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 43 152 44 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 48 611 49 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 578 48 71 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 49 152 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 72 71 74 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 578 77 72 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00068 73 595 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00067 74 79 73 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00066 578 74 70 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 101 62 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 578 55 58 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 58 56 62 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 61 473 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 578 528 57 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 62 64 61 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 57 70 62 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 578 164 54 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00057 56 54 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 578 340 56 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00055 52 71 53 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 53 349 52 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 52 586 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 578 620 50 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 50 577 51 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 578 59 63 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 63 60 64 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 107 528 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 578 340 107 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 66 614 65 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 65 67 66 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 66 473 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 578 107 47 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 47 44 46 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 46 45 60 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 45 42 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 42 595 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 578 155 42 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00037 578 39 40 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 39 80 578 578 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00035 578 614 349 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 141 38 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 38 604 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 578 40 38 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00031 578 75 80 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 34 528 20 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 578 34 138 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 20 604 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 578 176 10 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 578 566 18 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 18 611 19 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 578 614 8 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 8 138 7 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 7 19 59 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 578 10 9 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 9 611 11 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 578 604 16 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 16 349 17 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 27 528 12 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 578 27 28 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 12 566 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 578 595 6 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 6 17 5 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 5 51 55 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 578 595 611 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 578 65 1 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 1 261 24 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 24 22 578 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 15 51 578 578 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 14 349 13 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 578 15 14 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 578 13 2 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 2 11 4 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 4 28 3 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 3 53 22 578 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C625 10 578 5.489e-14
C624 11 578 5.436e-14
C622 13 578 5.826e-14
C620 15 578 1.662e-14
C618 17 578 5.566e-14
C616 19 578 5.226e-14
C612 22 578 7.271e-14
C610 24 578 2.773e-14
C609 25 578 6.05e-15
C607 27 578 1.8635e-14
C606 28 578 5.188e-14
C603 31 578 7.79e-15
C602 32 578 7.43e-15
C600 34 578 1.8635e-14
C597 37 578 7.43e-15
C596 38 578 1.8635e-14
C595 39 578 1.568e-14
C594 40 578 4.693e-14
C591 42 578 1.8635e-14
C589 44 578 5.326e-14
C588 45 578 5.876e-14
C585 48 578 1.8635e-14
C582 51 578 1.0199e-13
C581 52 578 4.11e-15
C580 53 578 6.152e-14
C579 54 578 1.677e-14
C578 55 578 5.1e-14
C577 56 578 4.738e-14
C574 59 578 5.945e-14
C573 60 578 1.067e-13
C571 62 578 2.9265e-14
C569 64 578 4.761e-14
C568 65 578 1.2107e-13
C567 66 578 4.11e-15
C566 67 578 4.997e-14
C565 68 578 4.11e-15
C564 69 578 1.853e-14
C563 70 578 7.468e-14
C562 71 578 1.541e-13
C559 74 578 2.445e-14
C558 75 578 1.0224e-13
C557 76 578 1.568e-14
C556 77 578 4.513e-14
C554 79 578 5.961e-14
C553 80 578 1.0734e-13
C552 81 578 1.8635e-14
C550 83 578 4.11e-15
C546 87 578 4.11e-15
C544 89 578 4.11e-15
C534 98 578 3.123e-14
C533 99 578 2.299e-14
C531 101 578 9.176e-14
C530 102 578 8.58e-15
C529 103 578 4.622e-14
C528 104 578 1.853e-14
C525 107 578 9.13e-14
C524 108 578 5.041e-14
C521 111 578 2.605e-14
C519 113 578 8.58e-15
C518 114 578 6.317e-14
C517 115 578 1.853e-14
C514 118 578 4.513e-14
C512 120 578 1.8635e-14
C509 123 578 7.56e-15
C508 124 578 2.596e-14
C507 125 578 7.76e-15
C506 126 578 4.835e-14
C504 128 578 5.387e-14
C503 129 578 2.16e-14
C502 130 578 1.8635e-14
C499 133 578 8.58e-15
C495 137 578 7.56e-15
C494 138 578 1.0967e-13
C491 141 578 1.0214e-13
C488 144 578 4.581e-14
C486 146 578 6.05e-15
C485 147 578 2.596e-14
C484 148 578 2.16e-14
C483 149 578 7.76e-15
C482 150 578 5.894e-14
C479 152 578 1.4772e-13
C478 153 578 1.8635e-14
C476 155 578 1.0282e-13
C475 156 578 6.122e-14
C474 157 578 1.853e-14
C473 158 578 4.11e-15
C472 159 578 7.479e-14
C471 160 578 1.27e-13
C470 161 578 4.11e-15
C468 163 578 2.299e-14
C467 164 578 1.3038e-13
C465 166 578 8.421e-14
C464 167 578 2.378e-14
C463 168 578 7.384e-14
C461 170 578 2.128e-14
C460 171 578 7.56e-15
C459 172 578 3.608e-14
C457 174 578 7.097e-14
C456 175 578 6.201e-14
C455 176 578 2.1142e-13
C453 178 578 2.299e-14
C452 179 578 4.11e-15
C451 180 578 6.578e-14
C450 181 578 7.532e-14
C448 183 578 2.378e-14
C446 185 578 3.608e-14
C445 186 578 7.56e-15
C443 188 578 2.128e-14
C442 189 578 4.112e-14
C441 190 578 7.43e-15
C440 191 578 2.455e-14
C439 192 578 1.3107e-13
C437 194 578 1.8635e-14
C436 195 578 5.953e-14
C435 196 578 9.133e-14
C434 197 578 1.8635e-14
C428 203 578 4.11e-15
C425 206 578 4.11e-15
C419 212 578 7.56e-15
C415 216 578 4.11e-15
C411 219 578 4.487e-14
C410 220 578 6.05e-15
C409 221 578 1.767e-14
C408 222 578 6.05e-15
C407 223 578 6.561e-14
C406 224 578 1.0793e-13
C405 225 578 9.158e-14
C404 226 578 7.523e-14
C403 227 578 1.853e-14
C401 229 578 1.8635e-14
C400 230 578 5.28e-14
C399 231 578 4.438e-14
C398 232 578 2.299e-14
C396 234 578 8.58e-15
C395 235 578 4.284e-14
C394 236 578 8.072e-14
C393 237 578 1.662e-14
C392 238 578 2.596e-14
C391 239 578 5.002e-14
C390 240 578 9.7e-15
C389 241 578 2.16e-14
C388 242 578 2.128e-14
C387 243 578 2.378e-14
C386 244 578 5.376e-14
C383 247 578 6.312e-14
C382 248 578 3.608e-14
C381 249 578 7.56e-15
C379 251 578 1.061e-13
C378 252 578 1.534e-13
C376 254 578 2.596e-14
C375 255 578 1.0305e-13
C374 256 578 9.7e-15
C373 257 578 2.16e-14
C371 259 578 7.43e-15
C369 261 578 1.0665e-13
C368 262 578 2.114e-13
C365 265 578 5.055e-14
C362 268 578 9.7e-15
C360 270 578 7.165e-14
C355 275 578 9.145e-14
C354 276 578 6.05e-15
C350 280 578 1.3368e-13
C344 286 578 7.877e-14
C342 288 578 6.05e-15
C340 290 578 5.043e-14
C339 291 578 6.05e-15
C337 293 578 1.0851e-13
C334 296 578 1.5036e-13
C333 297 578 4.11e-15
C330 299 578 5.107e-14
C329 300 578 2.445e-14
C327 302 578 2.605e-14
C323 306 578 2.596e-14
C322 307 578 2.16e-14
C321 308 578 1.8773e-13
C320 309 578 8.46e-14
C317 312 578 1.8635e-14
C314 315 578 5.535e-14
C313 316 578 2.605e-14
C312 317 578 2.455e-14
C310 319 578 6.1e-14
C309 320 578 5.492e-14
C308 321 578 7.361e-14
C307 322 578 1.767e-14
C304 325 578 1.767e-14
C301 328 578 1.853e-14
C298 330 578 2.596e-14
C297 331 578 5.125e-14
C296 332 578 2.16e-14
C295 333 578 9.7e-15
C294 334 578 8.086e-14
C293 335 578 6.05e-15
C292 336 578 5.283e-14
C291 337 578 1.8635e-14
C288 340 578 3.5983e-13
C287 341 578 6.072e-14
C286 342 578 2.455e-14
C285 343 578 8.1e-14
C284 344 578 5.779e-14
C283 345 578 6.066e-14
C282 346 578 6.05e-15
C281 347 578 1.1441e-13
C279 349 578 5.367e-13
C278 350 578 1.8635e-14
C276 352 578 5.495e-14
C275 353 578 7.42e-14
C274 354 578 6.05e-15
C273 355 578 1.0345e-13
C271 357 578 1.8635e-14
C270 358 578 2.596e-14
C269 359 578 9.7e-15
C268 360 578 2.16e-14
C267 361 578 1.0272e-13
C266 362 578 1.568e-14
C265 363 578 5.248e-14
C264 364 578 6.629e-14
C263 365 578 1.8635e-14
C262 366 578 1.318e-13
C261 367 578 1.568e-14
C260 368 578 5.395e-14
C259 369 578 9.7e-15
C257 371 578 1.0668e-13
C253 375 578 7.43e-15
C251 377 578 1.0173e-13
C248 380 578 7.56e-15
C244 384 578 4.11e-15
C243 385 578 1.7927e-13
C241 387 578 4.11e-15
C240 388 578 8.58e-15
C238 390 578 7.832e-14
C235 393 578 7.56e-15
C231 396 578 6.05e-15
C230 397 578 2.596e-14
C229 398 578 2.16e-14
C228 399 578 1.3174e-13
C226 401 578 1.8635e-14
C225 402 578 5.169e-14
C221 406 578 1.568e-14
C220 407 578 4.971e-14
C219 408 578 4.11e-15
C218 409 578 2.445e-14
C217 410 578 1.1694e-13
C216 411 578 9.277e-14
C215 412 578 1.1703e-13
C214 413 578 4.11e-15
C213 414 578 2.378e-14
C212 415 578 5.874e-14
C208 419 578 2.128e-14
C207 420 578 8.106e-14
C206 421 578 6.4e-14
C204 423 578 3.608e-14
C203 424 578 7.56e-15
C199 428 578 1.853e-14
C196 431 578 5.102e-14
C195 432 578 8.897e-14
C194 433 578 2.299e-14
C192 435 578 1.8635e-14
C191 436 578 4.558e-14
C189 438 578 4.11e-15
C188 439 578 9.206e-14
C187 440 578 2.378e-14
C184 443 578 2.128e-14
C183 444 578 7.56e-15
C181 446 578 3.608e-14
C179 448 578 4.0274e-13
C178 449 578 7.56e-15
C175 452 578 5.061e-14
C174 453 578 5.113e-14
C172 455 578 9.643e-14
C170 456 578 4.489e-14
C168 458 578 8.188e-14
C167 459 578 1.8635e-14
C166 460 578 5.233e-14
C165 461 578 1.0783e-13
C162 464 578 6.632e-14
C161 465 578 5.011e-14
C159 467 578 5.532e-14
C158 468 578 8.817e-14
C157 469 578 5.865e-14
C156 470 578 5.247e-14
C155 471 578 2.605e-14
C154 472 578 2.678e-13
C153 473 578 5.8288e-13
C152 474 578 2.605e-14
C150 476 578 1.8635e-14
C149 477 578 1.0692e-13
C148 478 578 6.56e-14
C146 480 578 4.363e-14
C145 481 578 1.568e-14
C144 482 578 9.642e-14
C143 483 578 5.972e-14
C141 485 578 5.232e-14
C140 486 578 2.378e-14
C139 487 578 2.128e-14
C137 489 578 3.608e-14
C135 491 578 7.56e-15
C134 492 578 1.2768e-13
C133 493 578 4.72e-14
C131 495 578 7.56e-15
C127 499 578 9.7e-15
C126 500 578 9.7e-15
C125 501 578 7.43e-15
C123 503 578 9.7e-15
C122 504 578 7.76e-15
C121 505 578 9.7e-15
C119 507 578 7.76e-15
C117 508 578 1.8635e-14
C115 510 578 4.6496e-13
C114 511 578 2.378e-14
C113 512 578 7.221e-14
C111 514 578 2.128e-14
C109 516 578 7.56e-15
C107 518 578 3.608e-14
C105 520 578 4.7208e-13
C104 521 578 4.891e-14
C103 522 578 2.596e-14
C102 523 578 5.486e-14
C100 525 578 2.16e-14
C98 527 578 4.11e-15
C97 528 578 7.56709e-13
C95 530 578 6.07e-14
C93 532 578 2.596e-14
C92 533 578 2.16e-14
C91 534 578 5.169e-14
C90 535 578 4.11e-15
C88 537 578 2.445e-14
C84 541 578 5.775e-14
C80 545 578 2.3093e-13
C79 546 578 4.11e-15
C78 547 578 2.596e-14
C77 548 578 1.219e-13
C76 549 578 6.445e-14
C74 551 578 2.16e-14
C71 554 578 2.596e-14
C70 555 578 4.11e-15
C68 557 578 2.16e-14
C67 558 578 2.596e-14
C66 559 578 5.913e-14
C64 561 578 2.16e-14
C62 563 578 4.11e-15
C61 564 578 1.2557e-13
C59 566 578 4.8009e-13
C58 567 578 1.8635e-14
C54 571 578 2.596e-14
C52 573 578 6.3875e-13
C51 574 578 5.937e-14
C49 576 578 2.16e-14
C48 577 578 6.1861e-13
C47 578 578 7.21657e-12
C46 579 578 3.139e-14
C45 580 578 1.8635e-14
C43 582 578 5.676e-14
C42 583 578 9.182e-14
C41 584 578 5.713e-14
C39 586 578 3.6947e-13
C38 587 578 5.979e-14
C36 589 578 5.025e-14
C35 590 578 7.912e-14
C34 591 578 2.605e-14
C33 592 578 5.892e-14
C32 593 578 6.152e-14
C31 594 578 1.0514e-13
C30 595 578 1.24632e-12
C28 597 578 2.455e-14
C26 599 578 6.073e-14
C25 600 578 6.547e-14
C24 601 578 1.853e-14
C21 604 578 1.19869e-12
C20 605 578 1.7998e-13
C19 606 578 8.018e-14
C18 607 578 1.8635e-14
C17 608 578 1.0517e-13
C16 609 578 1.853e-14
C14 611 578 1.05486e-12
C13 612 578 1.4686e-13
C12 613 578 1.8635e-14
C11 614 578 8.81409e-13
C10 615 578 2.596e-14
C9 616 578 5.001e-14
C8 617 578 9.7e-15
C7 618 578 2.16e-14
C6 619 578 7.929e-14
C5 620 578 9.40519e-13
C4 621 578 5.8358e-13
C3 622 578 7.47362e-12
C2 623 578 6.057e-14
.ends mul4b_cougar

