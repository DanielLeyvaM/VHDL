* Spice description of act5_cougar
* Spice driver version -1208783196
* Date ( dd/mm/yyyy hh:mm:ss ): 23/11/2020 at 13:04:07

* INTERF clk ctrl ctrl1 dh[0] dh[1] dh[2] dh[3] dm[0] dm[1] dm[2] dm[3] rst 
* INTERF uh[0] uh[1] uh[2] uh[3] um[0] um[1] um[2] um[3] vdd vss 


.subckt act5_cougar 1881 1111 187 364 309 188 463 1230 1148 1056 957 1845 831 761 647 465 1804 1653 1507 1394 1885 1803 
* NET 24 = not_maquina
* NET 26 = mbk_buf_not_maquina
* NET 30 = not_aux15
* NET 34 = mbk_buf_aux16
* NET 38 = a3_x2_8_sig
* NET 39 = no3_x1_8_sig
* NET 43 = cum_2_ins.sff_s
* NET 44 = cum_2_ins.y
* NET 45 = cum_2_ins.sff_m
* NET 48 = oa22_x2_4_sig
* NET 49 = cum_2_ins.u
* NET 50 = cum_2_ins.nckr
* NET 51 = cum_2_ins.ckr
* NET 53 = maquina
* NET 55 = maquina_ins.sff_s
* NET 57 = maquina_ins.y
* NET 59 = maquina_ins.sff_m
* NET 62 = maquina_ins.nckr
* NET 63 = maquina_ins.u
* NET 64 = maquina_ins.ckr
* NET 69 = cdm_0_ins.y
* NET 71 = cdm_0_ins.sff_m
* NET 73 = cdm_0_ins.sff_s
* NET 74 = cdm_0_ins.u
* NET 75 = cdm_0_ins.ckr
* NET 76 = cdm_0_ins.nckr
* NET 77 = no2_x1_6_sig
* NET 80 = mbk_buf_mbk_buf_maquina
* NET 83 = nxr2_x1_2_sig
* NET 85 = cum_1_ins.sff_s
* NET 86 = cum_1_ins.y
* NET 89 = cum_1_ins.sff_m
* NET 90 = cum_1_ins.nckr
* NET 91 = cum_1_ins.u
* NET 92 = cum_1_ins.ckr
* NET 93 = mbk_buf_maquina
* NET 96 = aux0
* NET 102 = nao2o22_x1_sig
* NET 104 = o3_x2_5_sig
* NET 112 = not_aux71
* NET 114 = noa22_x1_sig
* NET 117 = o3_x2_6_sig
* NET 118 = not_aux147
* NET 122 = not_aux58
* NET 125 = o2_x2_8_sig
* NET 130 = no2_x1_22_sig
* NET 131 = na2_x1_18_sig
* NET 134 = nao22_x1_6_sig
* NET 135 = oa2a22_x2_sig
* NET 139 = cum_3_ins.sff_s
* NET 140 = cum_3_ins.y
* NET 143 = cum_3_ins.sff_m
* NET 144 = oa22_x2_5_sig
* NET 145 = cum_3_ins.u
* NET 146 = cum_3_ins.ckr
* NET 147 = cum_3_ins.nckr
* NET 148 = na3_x1_13_sig
* NET 150 = na3_x1_12_sig
* NET 155 = na3_x1_14_sig
* NET 157 = na2_x1_11_sig
* NET 187 = ctrl1
* NET 188 = dh[2]
* NET 189 = cum[0]
* NET 192 = cum_0_ins.sff_s
* NET 193 = cum_0_ins.y
* NET 195 = cum_0_ins.sff_m
* NET 197 = cum_0_ins.u
* NET 198 = cum_0_ins.ckr
* NET 200 = na2_x1_16_sig
* NET 201 = cum_0_ins.nckr
* NET 202 = mbk_buf_aux0
* NET 203 = na3_x1_18_sig
* NET 204 = no2_x1_21_sig
* NET 208 = no3_x1_7_sig
* NET 211 = not_aux0
* NET 212 = an12_x1_2_sig
* NET 217 = cdm_3_ins.sff_s
* NET 218 = cdm_3_ins.y
* NET 219 = cdm_3_ins.u
* NET 221 = cdm_3_ins.sff_m
* NET 223 = aux16
* NET 224 = cdm_3_ins.nckr
* NET 225 = cdm_3_ins.ckr
* NET 226 = cum[1]
* NET 231 = na2_x1_10_sig
* NET 232 = na2_x1_15_sig
* NET 233 = nao22_x1_5_sig
* NET 234 = oa22_x2_3_sig
* NET 238 = not_aux70
* NET 241 = a4_x2_sig
* NET 242 = no2_x1_17_sig
* NET 244 = aux150
* NET 247 = oa22_x2_2_sig
* NET 248 = na2_x1_12_sig
* NET 250 = na3_x1_16_sig
* NET 251 = not_aux59
* NET 253 = no2_x1_19_sig
* NET 255 = on12_x1_4_sig
* NET 257 = cdm_1_ins.y
* NET 259 = cdm_1_ins.sff_m
* NET 260 = cdm_1_ins.sff_s
* NET 261 = na3_x1_15_sig
* NET 262 = cdm_1_ins.u
* NET 264 = cdm_1_ins.nckr
* NET 265 = cdm_1_ins.ckr
* NET 266 = no2_x1_18_sig
* NET 272 = stop_ins.u
* NET 273 = stop_ins.ckr
* NET 274 = stop_ins.nckr
* NET 276 = na2_x1_17_sig
* NET 278 = mbk_buf_not_aux0
* NET 279 = no2_x1_7_sig
* NET 286 = not_aux39
* NET 292 = not_aux17
* NET 302 = na2_x1_14_sig
* NET 306 = not_aux60
* NET 309 = dh[1]
* NET 310 = stop_ins.sff_s
* NET 313 = stop_ins.sff_m
* NET 315 = stop_ins.y
* NET 321 = ao22_x2_sig
* NET 325 = aux146
* NET 327 = a2_x2_2_sig
* NET 333 = not_aux61
* NET 336 = o3_x2_3_sig
* NET 345 = not_aux19
* NET 352 = aux64
* NET 354 = nao22_x1_4_sig
* NET 358 = no2_x1_20_sig
* NET 359 = na3_x1_17_sig
* NET 364 = dh[0]
* NET 367 = rtlalc_9_1_ins.sff_s
* NET 368 = rtlalc_9_1_ins.y
* NET 370 = rtlalc_9_1_ins.sff_m
* NET 371 = rtlalc_9_1_ins.u
* NET 373 = rtlalc_9_1_ins.ckr
* NET 374 = not_cum[0]
* NET 375 = rtlalc_9_1_ins.nckr
* NET 376 = not_cum[1]
* NET 378 = not_aux145
* NET 380 = inv_x2_2_sig
* NET 381 = not_aux1
* NET 383 = mbk_buf_not_aux1
* NET 386 = aux11
* NET 389 = not_aux42
* NET 390 = not_stop
* NET 391 = na4_x1_5_sig
* NET 392 = na2_x1_5_sig
* NET 393 = no2_x1_10_sig
* NET 397 = on12_x1_2_sig
* NET 399 = mbk_buf_not_aux15
* NET 400 = no2_x1_11_sig
* NET 402 = o3_x2_2_sig
* NET 407 = cdh[2]
* NET 409 = cdh_2_ins.sff_s
* NET 410 = cdh_2_ins.y
* NET 412 = cdh_2_ins.sff_m
* NET 414 = oa3ao322_x2_sig
* NET 415 = cdh_2_ins.nckr
* NET 416 = cdh_2_ins.u
* NET 417 = cdh_2_ins.ckr
* NET 418 = aux66
* NET 419 = not_cdm[2]
* NET 420 = inv_x2_4_sig
* NET 424 = o3_x2_4_sig
* NET 425 = a4_x2_4_sig
* NET 427 = cdm_2_ins.sff_s
* NET 428 = cdm_2_ins.y
* NET 430 = cdm_2_ins.sff_m
* NET 431 = na2_x1_13_sig
* NET 432 = cdm_2_ins.u
* NET 434 = cdm_2_ins.ckr
* NET 435 = cdm_2_ins.nckr
* NET 463 = dh[3]
* NET 465 = uh[3]
* NET 469 = rtlalc_9_2_ins.sff_s
* NET 470 = rtlalc_9_2_ins.y
* NET 471 = rtlalc_9_2_ins.sff_m
* NET 477 = rtlalc_9_2_ins.nckr
* NET 478 = rtlalc_9_2_ins.u
* NET 479 = rtlalc_9_2_ins.ckr
* NET 482 = cdh_1_ins.sff_s
* NET 484 = cdh_1_ins.y
* NET 485 = cdh_1_ins.sff_m
* NET 488 = cdh_1_ins.nckr
* NET 489 = cdh_1_ins.u
* NET 490 = cdh_1_ins.ckr
* NET 495 = cdh[1]
* NET 498 = o3_x2_sig
* NET 500 = nao22_x1_sig
* NET 501 = an12_x1_sig
* NET 508 = na4_x1_sig
* NET 511 = cum[2]
* NET 513 = no2_x1_4_sig
* NET 514 = no2_x1_3_sig
* NET 517 = na4_x1_2_sig
* NET 520 = a2_x2_sig
* NET 524 = na4_x1_4_sig
* NET 526 = no3_x1_4_sig
* NET 527 = no3_x1_3_sig
* NET 531 = no4_x1_5_sig
* NET 532 = no3_x1_sig
* NET 533 = na2_x1_4_sig
* NET 534 = stop
* NET 535 = no3_x1_2_sig
* NET 537 = na2_x1_3_sig
* NET 544 = not_aux47
* NET 552 = cuh_2_ins.sff_m
* NET 553 = cuh_2_ins.y
* NET 554 = cuh_2_ins.sff_s
* NET 556 = cuh_2_ins.u
* NET 557 = cuh_2_ins.ckr
* NET 558 = cuh_2_ins.nckr
* NET 560 = rtlalc_9[2]
* NET 561 = rtlalc_9[1]
* NET 563 = na2_x1_24_sig
* NET 564 = na3_x1_25_sig
* NET 565 = not_aux25
* NET 566 = aux139
* NET 567 = na3_x1_24_sig
* NET 569 = no2_x1_35_sig
* NET 572 = no3_x1_14_sig
* NET 573 = no2_x1_34_sig
* NET 575 = oa2a22_x2_3_sig
* NET 576 = not_rtlalc_9[2]
* NET 579 = aux24
* NET 581 = a2_x2_7_sig
* NET 583 = not_cdh[2]
* NET 584 = not_cdh[1]
* NET 588 = mbk_buf_not_aux17
* NET 589 = no4_x1_6_sig
* NET 590 = no2_x1_12_sig
* NET 591 = na4_x1_6_sig
* NET 592 = na2_x1_6_sig
* NET 595 = cdh_3_ins.sff_s
* NET 596 = nao22_x1_2_sig
* NET 597 = cdh_3_ins.y
* NET 600 = cdh_3_ins.sff_m
* NET 601 = cdh_3_ins.u
* NET 602 = cdh_3_ins.nckr
* NET 603 = cdh_3_ins.ckr
* NET 604 = cdm[3]
* NET 606 = no3_x1_5_sig
* NET 608 = o4_x2_2_sig
* NET 615 = aux48
* NET 616 = na3_x1_10_sig
* NET 617 = na3_x1_9_sig
* NET 618 = not_aux56
* NET 619 = not_aux49
* NET 622 = o2_x2_6_sig
* NET 623 = on12_x1_3_sig
* NET 647 = uh[2]
* NET 652 = rtlalc_9_0_ins.sff_m
* NET 653 = rtlalc_9_0_ins.sff_s
* NET 655 = rtlalc_9_0_ins.y
* NET 656 = rtlalc_9_0_ins.u
* NET 658 = rtlalc_9_0_ins.ckr
* NET 661 = rtlalc_9[0]
* NET 662 = rtlalc_9_0_ins.nckr
* NET 664 = no2_x1_33_sig
* NET 665 = no3_x1_12_sig
* NET 666 = rtlalc_9_3_ins.y
* NET 667 = rtlalc_9_3_ins.sff_s
* NET 669 = rtlalc_9_3_ins.u
* NET 671 = rtlalc_9_3_ins.sff_m
* NET 673 = rtlalc_9[3]
* NET 674 = rtlalc_9_3_ins.nckr
* NET 675 = rtlalc_9_3_ins.ckr
* NET 677 = no2_x1_36_sig
* NET 678 = no3_x1_15_sig
* NET 682 = a2_x2_11_sig
* NET 684 = cdh[3]
* NET 685 = not_cdh[3]
* NET 687 = o2_x2_3_sig
* NET 688 = an12_x1_4_sig
* NET 690 = no2_x1_9_sig
* NET 691 = mbk_buf_aux21
* NET 695 = not_aux10
* NET 697 = a4_x2_3_sig
* NET 701 = a3_x2_4_sig
* NET 703 = aux21
* NET 707 = not_aux43
* NET 710 = cdm[0]
* NET 711 = o2_x2_5_sig
* NET 716 = not_aux54
* NET 719 = na2_x1_8_sig
* NET 720 = no2_x1_14_sig
* NET 726 = na3_x1_7_sig
* NET 727 = o2_x2_4_sig
* NET 728 = na3_x1_8_sig
* NET 732 = cuh_1_ins.y
* NET 734 = cuh_1_ins.sff_m
* NET 735 = cuh_1_ins.sff_s
* NET 738 = na3_x1_6_sig
* NET 740 = cuh_1_ins.u
* NET 741 = cuh_1_ins.ckr
* NET 742 = cuh_1_ins.nckr
* NET 751 = na2_x1_28_sig
* NET 753 = na2_x1_29_sig
* NET 755 = na2_x1_27_sig
* NET 757 = mbk_buf_not_aux19
* NET 759 = no2_x1_15_sig
* NET 761 = uh[1]
* NET 762 = rtlalc_10[2]
* NET 763 = rtlalc_10_2_ins.ckr
* NET 764 = rtlalc_10_2_ins.nckr
* NET 765 = rtlalc_10_2_ins.sff_m
* NET 767 = rtlalc_10_2_ins.y
* NET 769 = rtlalc_10_2_ins.sff_s
* NET 770 = rtlalc_10_2_ins.u
* NET 774 = o2_x2_14_sig
* NET 777 = no3_x1_13_sig
* NET 781 = a3_x2_14_sig
* NET 782 = rtlalc_10_1_ins.ckr
* NET 786 = rtlalc_10_1_ins.nckr
* NET 787 = rtlalc_10_1_ins.sff_m
* NET 788 = rtlalc_10_1_ins.sff_s
* NET 789 = rtlalc_10_1_ins.y
* NET 793 = rtlalc_10_1_ins.u
* NET 796 = o2_x2_13_sig
* NET 799 = a3_x2_13_sig
* NET 804 = not_cuh[1]
* NET 805 = o2_x2_7_sig
* NET 806 = no4_x1_7_sig
* NET 810 = no2_x1_16_sig
* NET 812 = cdm[1]
* NET 813 = not_cuh[0]
* NET 815 = no2_x1_8_sig
* NET 821 = inv_x2_3_sig
* NET 822 = o2_x2_sig
* NET 824 = no4_x1_4_sig
* NET 828 = cuh[2]
* NET 831 = uh[0]
* NET 834 = aux140
* NET 838 = na3_x1_27_sig
* NET 839 = na3_x1_26_sig
* NET 841 = rtlalc_10[0]
* NET 842 = rtlalc_10_0_ins.y
* NET 843 = rtlalc_10_0_ins.sff_s
* NET 845 = na2_x1_25_sig
* NET 846 = rtlalc_10_0_ins.u
* NET 848 = rtlalc_10_0_ins.sff_m
* NET 850 = rtlalc_10_0_ins.ckr
* NET 853 = rtlalc_10_0_ins.nckr
* NET 854 = not_cdm[3]
* NET 856 = na2_x1_37_sig
* NET 857 = no3_x1_16_sig
* NET 860 = rtlalc_10_3_ins.y
* NET 862 = rtlalc_10_3_ins.sff_m
* NET 863 = rtlalc_10_3_ins.sff_s
* NET 864 = rtlalc_10_3_ins.u
* NET 866 = rtlalc_10_3_ins.ckr
* NET 867 = not_aux138
* NET 869 = rtlalc_10_3_ins.nckr
* NET 870 = na2_x1_31_sig
* NET 872 = na3_x1_28_sig
* NET 874 = na2_x1_30_sig
* NET 878 = a3_x2_5_sig
* NET 879 = aux63
* NET 886 = a4_x2_2_sig
* NET 889 = aux57
* NET 891 = not_cdm[0]
* NET 892 = cuh[1]
* NET 894 = not_aux14
* NET 897 = na2_x1_9_sig
* NET 898 = na3_x1_11_sig
* NET 903 = cuh_3_ins.y
* NET 904 = cuh_3_ins.sff_s
* NET 906 = na4_x1_8_sig
* NET 907 = cuh_3_ins.u
* NET 908 = cuh_3_ins.ckr
* NET 909 = cuh_3_ins.sff_m
* NET 911 = cuh_3_ins.nckr
* NET 912 = oa22_x2_sig
* NET 914 = nxr2_x1_3_sig
* NET 915 = nao22_x1_3_sig
* NET 918 = cuh[3]
* NET 931 = rtlalc_10[1]
* NET 957 = dm[3]
* NET 962 = rtlalc_11[3]
* NET 964 = rtlalc_11_3_ins.sff_s
* NET 967 = rtlalc_11_3_ins.y
* NET 969 = rtlalc_11_3_ins.sff_m
* NET 970 = rtlalc_11_3_ins.u
* NET 971 = rtlalc_11_3_ins.nckr
* NET 972 = rtlalc_11_3_ins.ckr
* NET 974 = na3_x1_32_sig
* NET 975 = na2_x1_35_sig
* NET 977 = aux141
* NET 978 = na3_x1_31_sig
* NET 981 = o3_x2_8_sig
* NET 982 = an12_x1_5_sig
* NET 986 = na2_x1_36_sig
* NET 988 = rtlalc_11_2_ins.sff_s
* NET 990 = rtlalc_11_2_ins.y
* NET 991 = rtlalc_11_2_ins.u
* NET 992 = rtlalc_11_2_ins.sff_m
* NET 996 = rtlalc_11_2_ins.nckr
* NET 997 = rtlalc_11_2_ins.ckr
* NET 999 = na2_x1_33_sig
* NET 1000 = na3_x1_30_sig
* NET 1003 = na2_x1_34_sig
* NET 1006 = a2_x2_4_sig
* NET 1008 = a3_x2_6_sig
* NET 1012 = a2_x2_6_sig
* NET 1013 = a2_x2_5_sig
* NET 1015 = cum[3]
* NET 1016 = not_cum[3]
* NET 1020 = na3_x1_4_sig
* NET 1023 = na4_x1_3_sig
* NET 1026 = a2_x2_3_sig
* NET 1027 = na3_x1_3_sig
* NET 1029 = not_cuh[2]
* NET 1030 = na2_x1_2_sig
* NET 1031 = not_aux21
* NET 1033 = a3_x2_3_sig
* NET 1034 = not_cdm[1]
* NET 1035 = cdm[2]
* NET 1036 = not_aux149
* NET 1040 = rtlalc_11_1_ins.sff_s
* NET 1041 = rtlalc_11_1_ins.y
* NET 1042 = rtlalc_11_1_ins.u
* NET 1043 = rtlalc_11_1_ins.sff_m
* NET 1046 = rtlalc_11_1_ins.ckr
* NET 1047 = rtlalc_11_1_ins.nckr
* NET 1049 = a3_x2_16_sig
* NET 1051 = o2_x2_16_sig
* NET 1052 = o3_x2_12_sig
* NET 1056 = dm[2]
* NET 1059 = na3_x1_29_sig
* NET 1064 = na3_x1_37_sig
* NET 1065 = na3_x1_36_sig
* NET 1067 = aux144
* NET 1068 = not_cum[2]
* NET 1069 = na2_x1_42_sig
* NET 1072 = rtlalc_10[3]
* NET 1073 = o3_x2_10_sig
* NET 1074 = no2_x1_37_sig
* NET 1075 = o2_x2_17_sig
* NET 1079 = mdh_3_ins.y
* NET 1080 = mdh_3_ins.sff_s
* NET 1081 = mdh_3_ins.u
* NET 1084 = mdh_3_ins.sff_m
* NET 1085 = mdh_3_ins.ckr
* NET 1086 = mdh_3_ins.nckr
* NET 1087 = rtlalc_11[2]
* NET 1088 = o3_x2_13_sig
* NET 1089 = no2_x1_38_sig
* NET 1092 = cdh_0_ins.sff_s
* NET 1093 = cdh_0_ins.y
* NET 1095 = cdh_0_ins.sff_m
* NET 1097 = na3_x1_2_sig
* NET 1098 = cdh_0_ins.nckr
* NET 1099 = cdh_0_ins.u
* NET 1100 = cdh_0_ins.ckr
* NET 1101 = cdh[0]
* NET 1103 = o2_x2_2_sig
* NET 1104 = not_aux23
* NET 1105 = na4_x1_7_sig
* NET 1109 = ao22_x2_2_sig
* NET 1111 = ctrl
* NET 1148 = dm[1]
* NET 1149 = rtlalc_11[1]
* NET 1150 = not_maquina1
* NET 1151 = na2_x1_26_sig
* NET 1154 = na2_x1_40_sig
* NET 1155 = aux143
* NET 1156 = na3_x1_34_sig
* NET 1157 = na3_x1_35_sig
* NET 1159 = rtlalc_12_1_ins.sff_s
* NET 1160 = rtlalc_12_1_ins.y
* NET 1162 = rtlalc_12_1_ins.sff_m
* NET 1164 = na2_x1_39_sig
* NET 1165 = rtlalc_12_1_ins.nckr
* NET 1166 = rtlalc_12_1_ins.u
* NET 1167 = rtlalc_12_1_ins.ckr
* NET 1169 = rtlalc_12[2]
* NET 1170 = rtlalc_12_2_ins.y
* NET 1172 = rtlalc_12_2_ins.sff_s
* NET 1175 = na2_x1_41_sig
* NET 1176 = rtlalc_12_2_ins.u
* NET 1178 = rtlalc_12_2_ins.sff_m
* NET 1179 = rtlalc_12_2_ins.ckr
* NET 1181 = o2_x2_12_sig
* NET 1182 = rtlalc_12_2_ins.nckr
* NET 1184 = na2_x1_21_sig
* NET 1185 = na3_x1_21_sig
* NET 1187 = oa22_x2_7_sig
* NET 1188 = nao22_x1_8_sig
* NET 1193 = no3_x1_11_sig
* NET 1194 = not_muh[3]
* NET 1195 = not_mdh[3]
* NET 1197 = mdm_1_ins.y
* NET 1198 = mdm_1_ins.sff_s
* NET 1200 = mdm_1_ins.u
* NET 1202 = mdm_1_ins.sff_m
* NET 1203 = mdm_1_ins.ckr
* NET 1205 = mdm_1_ins.nckr
* NET 1207 = not_aux44
* NET 1208 = mbk_buf_not_aux47
* NET 1212 = a3_x2_7_sig
* NET 1213 = no3_x1_6_sig
* NET 1215 = no2_x1_13_sig
* NET 1216 = na2_x1_7_sig
* NET 1217 = not_aux38
* NET 1218 = cuh[0]
* NET 1221 = cuh_0_ins.y
* NET 1223 = cuh_0_ins.sff_m
* NET 1224 = cuh_0_ins.sff_s
* NET 1225 = na3_x1_5_sig
* NET 1227 = cuh_0_ins.nckr
* NET 1228 = cuh_0_ins.u
* NET 1229 = cuh_0_ins.ckr
* NET 1230 = dm[0]
* NET 1235 = rtlalc_11_0_ins.u
* NET 1236 = rtlalc_11_0_ins.ckr
* NET 1239 = rtlalc_11_0_ins.nckr
* NET 1240 = o2_x2_15_sig
* NET 1241 = na2_x1_32_sig
* NET 1244 = a3_x2_15_sig
* NET 1245 = rtlalc_11[0]
* NET 1247 = o3_x2_11_sig
* NET 1249 = an12_x1_6_sig
* NET 1252 = o3_x2_9_sig
* NET 1258 = rtlalc_12_3_ins.u
* NET 1262 = rtlalc_12_3_ins.ckr
* NET 1263 = rtlalc_12_3_ins.nckr
* NET 1264 = na2_x1_43_sig
* NET 1267 = a3_x2_17_sig
* NET 1268 = o2_x2_18_sig
* NET 1271 = o3_x2_14_sig
* NET 1274 = not_aux78
* NET 1281 = no2_x1_24_sig
* NET 1283 = na3_x1_19_sig
* NET 1287 = oa2a22_x2_2_sig
* NET 1288 = na2_x1_23_sig
* NET 1295 = no4_x1_8_sig
* NET 1298 = inv_x2_sig
* NET 1303 = mum_0_ins.u
* NET 1304 = mum_0_ins.ckr
* NET 1306 = nxr2_x1_sig
* NET 1308 = mum_0_ins.nckr
* NET 1313 = no2_x1_5_sig
* NET 1314 = maquina1_ins.u
* NET 1315 = maquina1_ins.ckr
* NET 1316 = maquina1_ins.nckr
* NET 1319 = rtlalc_11_0_ins.sff_s
* NET 1321 = rtlalc_11_0_ins.y
* NET 1322 = rtlalc_11_0_ins.sff_m
* NET 1334 = rtlalc_12_3_ins.sff_s
* NET 1335 = rtlalc_12_3_ins.y
* NET 1336 = rtlalc_12_3_ins.sff_m
* NET 1353 = a2_x2_8_sig
* NET 1354 = no3_x1_9_sig
* NET 1355 = a4_x2_5_sig
* NET 1361 = mum_0_ins.sff_s
* NET 1363 = mum_0_ins.y
* NET 1364 = mum_0_ins.sff_m
* NET 1367 = maquina1_ins.sff_s
* NET 1369 = maquina1_ins.y
* NET 1370 = maquina1_ins.sff_m
* NET 1374 = rtlalc_12_0_ins.sff_s
* NET 1375 = rtlalc_12_0_ins.y
* NET 1376 = rtlalc_12_0_ins.u
* NET 1378 = rtlalc_12_0_ins.sff_m
* NET 1380 = rtlalc_12_0_ins.ckr
* NET 1381 = rtlalc_12_0_ins.nckr
* NET 1382 = na2_x1_38_sig
* NET 1384 = na3_x1_33_sig
* NET 1385 = maquina1
* NET 1387 = nao22_x1_12_sig
* NET 1388 = aux142
* NET 1390 = on12_x1_5_sig
* NET 1391 = rtlalc_12[3]
* NET 1394 = um[3]
* NET 1395 = no3_x1_10_sig
* NET 1399 = mdh[3]
* NET 1405 = nao22_x1_7_sig
* NET 1406 = na3_x1_20_sig
* NET 1407 = na3_x1_sig
* NET 1408 = not_aux104
* NET 1410 = a3_x2_2_sig
* NET 1411 = not_mdh[2]
* NET 1416 = no4_x1_2_sig
* NET 1417 = mdh[2]
* NET 1419 = mdh_2_ins.y
* NET 1420 = mdh_2_ins.sff_s
* NET 1421 = oa22_x2_6_sig
* NET 1422 = mdh_2_ins.ckr
* NET 1423 = mdh_2_ins.u
* NET 1425 = mdh_2_ins.sff_m
* NET 1427 = mdh_2_ins.nckr
* NET 1432 = no2_x1_31_sig
* NET 1433 = not_mdm[2]
* NET 1436 = not_aux133
* NET 1441 = not_aux107
* NET 1443 = nao2o22_x1_3_sig
* NET 1444 = no4_x1_9_sig
* NET 1448 = not_aux134
* NET 1450 = mdm_2_ins.sff_s
* NET 1451 = mdm_2_ins.y
* NET 1453 = mdm_2_ins.sff_m
* NET 1454 = oa22_x2_9_sig
* NET 1455 = mdm_2_ins.u
* NET 1457 = mdm_2_ins.nckr
* NET 1458 = mdm_2_ins.ckr
* NET 1469 = inv_x2_6_sig
* NET 1470 = no2_x1_26_sig
* NET 1480 = na2_x1_20_sig
* NET 1482 = no2_x1_sig
* NET 1507 = um[2]
* NET 1508 = muh_1_ins.sff_s
* NET 1509 = muh_1_ins.sff_m
* NET 1510 = muh_1_ins.y
* NET 1511 = muh_1_ins.ckr
* NET 1512 = muh_1_ins.u
* NET 1513 = oa2ao222_x2_3_sig
* NET 1517 = muh_1_ins.nckr
* NET 1522 = not_aux118
* NET 1524 = not_aux96
* NET 1527 = no4_x1_3_sig
* NET 1533 = no2_x1_2_sig
* NET 1534 = not_mdh[0]
* NET 1535 = na2_x1_sig
* NET 1540 = not_aux73
* NET 1548 = not_aux88
* NET 1551 = not_mdm[3]
* NET 1553 = not_aux148
* NET 1557 = no2_x1_32_sig
* NET 1559 = noa22_x1_3_sig
* NET 1561 = mdm[2]
* NET 1563 = not_aux116
* NET 1567 = not_aux132
* NET 1570 = mdm_3_ins.sff_s
* NET 1571 = mdm_3_ins.sff_m
* NET 1573 = mdm_3_ins.u
* NET 1574 = nao2o22_x1_4_sig
* NET 1575 = mdm_3_ins.y
* NET 1576 = mdm_3_ins.ckr
* NET 1579 = mdm_3_ins.nckr
* NET 1584 = mum_2_ins.sff_s
* NET 1586 = mum_2_ins.sff_m
* NET 1587 = mum_2_ins.ckr
* NET 1589 = mum_2_ins.y
* NET 1591 = mum_2_ins.u
* NET 1592 = nao22_x1_10_sig
* NET 1593 = mum_2_ins.nckr
* NET 1595 = rtlalc_12[0]
* NET 1596 = rtlalc_12[1]
* NET 1601 = nxr2_x1_4_sig
* NET 1604 = no2_x1_27_sig
* NET 1610 = o4_x2_sig
* NET 1611 = not_aux119
* NET 1613 = not_muh[1]
* NET 1615 = on12_x1_sig
* NET 1616 = a3_x2_sig
* NET 1619 = not_aux81
* NET 1620 = mdm[3]
* NET 1623 = na2_x1_19_sig
* NET 1624 = not_aux92
* NET 1626 = not_aux85
* NET 1627 = no4_x1_sig
* NET 1629 = inv_x2_7_sig
* NET 1630 = not_aux113
* NET 1634 = na3_x1_22_sig
* NET 1635 = o2_x2_10_sig
* NET 1639 = xr2_x1_3_sig
* NET 1641 = na3_x1_23_sig
* NET 1642 = mdm[0]
* NET 1644 = mdm_0_ins.sff_s
* NET 1645 = mdm_0_ins.y
* NET 1646 = mdm_0_ins.sff_m
* NET 1648 = nao22_x1_9_sig
* NET 1649 = mdm_0_ins.u
* NET 1651 = mdm_0_ins.ckr
* NET 1652 = mdm_0_ins.nckr
* NET 1653 = um[1]
* NET 1685 = muh_0_ins.sff_s
* NET 1687 = muh_0_ins.y
* NET 1688 = muh_0_ins.u
* NET 1690 = muh_0_ins.sff_m
* NET 1693 = muh_0_ins.ckr
* NET 1694 = muh_0_ins.nckr
* NET 1696 = a3_x2_10_sig
* NET 1700 = oa22_x2_8_sig
* NET 1702 = not_aux127
* NET 1703 = mdm[1]
* NET 1712 = a4_x2_6_sig
* NET 1713 = a3_x2_11_sig
* NET 1714 = no2_x1_30_sig
* NET 1715 = not_aux129
* NET 1719 = muh[3]
* NET 1722 = muh_3_ins.y
* NET 1724 = muh_3_ins.sff_m
* NET 1725 = muh_3_ins.sff_s
* NET 1728 = oa2ao222_x2_5_sig
* NET 1729 = muh_3_ins.u
* NET 1730 = muh_3_ins.ckr
* NET 1732 = not_aux111
* NET 1733 = nao2o22_x1_2_sig
* NET 1734 = muh_3_ins.nckr
* NET 1736 = not_mdh[1]
* NET 1737 = aux82
* NET 1740 = mdh_0_ins.y
* NET 1742 = mdh_0_ins.sff_s
* NET 1743 = mdh_0_ins.ckr
* NET 1744 = mdh_0_ins.u
* NET 1745 = mdh_0_ins.sff_m
* NET 1748 = mdh_0_ins.nckr
* NET 1749 = oa2ao222_x2_sig
* NET 1750 = an12_x1_3_sig
* NET 1751 = inv_x2_5_sig
* NET 1752 = mdh[0]
* NET 1756 = no2_x1_23_sig
* NET 1757 = noa22_x1_2_sig
* NET 1758 = a3_x2_9_sig
* NET 1763 = mdh[1]
* NET 1765 = mdh_1_ins.y
* NET 1767 = mdh_1_ins.sff_m
* NET 1768 = mdh_1_ins.sff_s
* NET 1770 = oa2ao222_x2_2_sig
* NET 1772 = mdh_1_ins.u
* NET 1773 = mdh_1_ins.ckr
* NET 1774 = mdh_1_ins.nckr
* NET 1778 = o3_x2_7_sig
* NET 1779 = not_mum[3]
* NET 1783 = not_rst
* NET 1787 = a3_x2_12_sig
* NET 1788 = nao22_x1_11_sig
* NET 1792 = mum[2]
* NET 1797 = xr2_x1_sig
* NET 1799 = not_aux137
* NET 1803 = vss
* NET 1804 = um[0]
* NET 1806 = muh[1]
* NET 1809 = xr2_x1_2_sig
* NET 1812 = a2_x2_9_sig
* NET 1813 = a2_x2_10_sig
* NET 1814 = no2_x1_28_sig
* NET 1818 = na2_x1_22_sig
* NET 1820 = no2_x1_29_sig
* NET 1822 = muh_2_ins.sff_s
* NET 1823 = muh_2_ins.y
* NET 1824 = oa2ao222_x2_4_sig
* NET 1826 = muh_2_ins.u
* NET 1828 = muh_2_ins.sff_m
* NET 1829 = muh_2_ins.nckr
* NET 1830 = muh_2_ins.ckr
* NET 1831 = not_muh[0]
* NET 1832 = o2_x2_9_sig
* NET 1833 = not_aux117
* NET 1836 = not_muh[2]
* NET 1837 = muh[2]
* NET 1840 = not_mdm[1]
* NET 1842 = muh[0]
* NET 1843 = not_mum[1]
* NET 1845 = rst
* NET 1846 = not_aux72
* NET 1849 = no2_x1_25_sig
* NET 1850 = not_mum[2]
* NET 1853 = not_aux105
* NET 1855 = not_aux131
* NET 1856 = not_aux130
* NET 1857 = o2_x2_11_sig
* NET 1858 = not_aux135
* NET 1861 = mum[1]
* NET 1863 = mum_1_ins.sff_s
* NET 1864 = mum_1_ins.y
* NET 1867 = mum_1_ins.sff_m
* NET 1868 = not_mum[0]
* NET 1869 = nao2o22_x1_5_sig
* NET 1870 = mum_1_ins.u
* NET 1871 = mum_1_ins.nckr
* NET 1872 = mum_1_ins.ckr
* NET 1873 = mum[0]
* NET 1875 = mum[3]
* NET 1876 = mum_3_ins.sff_s
* NET 1877 = mum_3_ins.y
* NET 1879 = mum_3_ins.sff_m
* NET 1880 = oa22_x2_10_sig
* NET 1881 = clk
* NET 1883 = mum_3_ins.u
* NET 1884 = mum_3_ins.ckr
* NET 1885 = vdd
* NET 1886 = mum_3_ins.nckr
Mtr_03768 1862 1861 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03767 1863 1872 1862 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03766 1864 1871 1863 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03765 1867 1871 1866 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03764 1866 1864 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03763 1865 1872 1867 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03762 1871 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03761 1885 1871 1872 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03760 1870 1869 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03759 1885 1870 1865 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03758 1885 1863 1861 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03757 1861 1863 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03756 1864 1867 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03755 1874 1875 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03754 1876 1884 1874 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03753 1877 1886 1876 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03752 1879 1886 1878 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03751 1878 1877 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03750 1882 1884 1879 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03749 1886 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03748 1885 1886 1884 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03747 1883 1880 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03746 1885 1883 1882 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03745 1885 1876 1875 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03744 1875 1876 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03743 1877 1879 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03742 1855 1856 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03741 1885 1873 1855 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03740 1844 1843 1847 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03739 1885 1845 1844 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03738 1858 1847 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03737 1852 1856 1854 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03736 1885 1853 1852 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03735 1857 1854 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03734 1869 1868 1860 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03733 1860 1857 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03732 1859 1858 1869 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03731 1885 1873 1859 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03730 1856 1851 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03729 1885 1850 1851 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03728 1851 1875 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03727 1868 1873 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03726 1848 1846 1849 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03725 1885 1845 1848 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03724 1838 1861 1839 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03723 1885 1845 1838 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03722 1853 1839 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03721 1834 1833 1835 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03720 1885 1845 1834 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03719 1832 1835 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03718 1836 1837 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03717 1843 1861 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03716 1805 1837 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03715 1885 1806 1808 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03714 1809 1805 1807 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03713 1807 1806 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03712 1807 1808 1809 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03711 1885 1837 1807 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03710 1818 1833 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03709 1885 1840 1818 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03708 1831 1842 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03707 1846 1841 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03706 1885 1840 1841 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03705 1841 1842 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03704 1813 1810 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03703 1885 1842 1810 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03702 1810 1809 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03701 1821 1837 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03700 1822 1830 1821 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03699 1823 1829 1822 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03698 1828 1829 1827 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03697 1827 1823 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03696 1825 1830 1828 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03695 1829 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03694 1885 1829 1830 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03693 1826 1824 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03692 1885 1826 1825 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03691 1885 1822 1837 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03690 1837 1822 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03689 1823 1828 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03688 1819 1836 1820 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03687 1885 1845 1819 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03686 1824 1815 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03685 1817 1812 1816 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03684 1817 1820 1885 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03683 1885 1818 1817 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03682 1816 1813 1815 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03681 1815 1814 1817 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03680 1812 1811 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03679 1885 1831 1811 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03678 1811 1837 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03677 1850 1792 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03676 1885 1797 1799 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03675 1799 1798 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03674 1885 1845 1798 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03673 1794 1792 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03672 1885 1861 1801 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03671 1797 1794 1683 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03670 1683 1861 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03669 1683 1801 1797 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03668 1885 1792 1683 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03667 1885 1790 1880 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03666 1682 1787 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03665 1682 1788 1790 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03664 1790 1873 1682 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03663 1673 1846 1756 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03662 1885 1845 1673 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03661 1885 1778 1788 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03660 1681 1779 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03659 1788 1799 1681 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03658 1779 1875 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03657 1885 1868 1786 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03656 1787 1786 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03655 1885 1783 1786 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03654 1786 1875 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03653 1885 1858 1680 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03652 1680 1875 1679 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03651 1679 1850 1776 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03650 1778 1776 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03649 1736 1763 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03648 1770 1760 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03647 1675 1758 1674 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03646 1675 1849 1885 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03645 1885 1763 1675 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03644 1674 1757 1760 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03643 1760 1846 1675 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03642 1749 1753 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03641 1671 1751 1672 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03640 1671 1756 1885 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03639 1885 1752 1671 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03638 1672 1750 1753 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03637 1753 1846 1671 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03636 1676 1763 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03635 1768 1773 1676 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03634 1765 1774 1768 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03633 1767 1774 1677 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03632 1677 1765 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03631 1678 1773 1767 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03630 1774 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03629 1885 1774 1773 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03628 1772 1770 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03627 1885 1772 1678 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03626 1885 1768 1763 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03625 1763 1768 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03624 1765 1767 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03623 1738 1737 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03622 1885 1738 1667 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03621 1667 1752 1750 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03620 1659 1715 1714 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03619 1885 1845 1659 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03618 1733 1831 1666 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03617 1666 1832 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03616 1665 1842 1733 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03615 1885 1732 1665 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03614 1885 1840 1707 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03613 1715 1707 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03612 1885 1833 1707 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03611 1707 1842 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03610 1662 1719 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03609 1725 1730 1662 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03608 1722 1734 1725 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03607 1724 1734 1663 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03606 1663 1722 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03605 1664 1730 1724 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03604 1734 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03603 1885 1734 1730 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03602 1729 1728 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03601 1885 1729 1664 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03600 1885 1725 1719 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03599 1719 1725 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03598 1722 1724 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03597 1728 1716 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03596 1661 1713 1660 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03595 1661 1714 1885 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03594 1885 1719 1661 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03593 1660 1712 1716 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03592 1716 1715 1661 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03591 1885 1705 1700 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03590 1658 1696 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03589 1658 1733 1705 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03588 1705 1840 1658 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03587 1657 1703 1814 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03586 1885 1702 1657 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03585 1669 1752 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03584 1742 1743 1669 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03583 1740 1748 1742 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03582 1745 1748 1668 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03581 1668 1740 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03580 1670 1743 1745 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03579 1748 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03578 1885 1748 1743 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03577 1744 1749 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03576 1885 1744 1670 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03575 1885 1742 1752 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03574 1752 1742 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03573 1740 1745 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03572 1885 1703 1699 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03571 1696 1699 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03570 1885 1783 1699 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03569 1699 1842 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03568 1654 1842 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03567 1685 1693 1654 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03566 1687 1694 1685 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03565 1690 1694 1656 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03564 1656 1687 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03563 1655 1693 1690 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03562 1694 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03561 1885 1694 1693 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03560 1688 1700 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03559 1885 1688 1655 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03558 1885 1685 1842 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03557 1842 1685 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03556 1687 1690 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03555 1885 1855 1634 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03554 1634 1642 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03553 1634 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03552 1637 1642 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03551 1885 1861 1640 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03550 1639 1637 1638 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03549 1638 1861 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03548 1638 1640 1639 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03547 1885 1642 1638 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03546 1643 1642 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03545 1644 1651 1643 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03544 1645 1652 1644 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03543 1646 1652 1647 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03542 1647 1645 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03541 1650 1651 1646 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03540 1652 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03539 1885 1652 1651 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03538 1649 1648 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03537 1885 1649 1650 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03536 1885 1644 1642 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03535 1642 1644 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03534 1645 1646 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03533 1632 1855 1633 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03532 1885 1845 1632 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03531 1635 1633 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03530 1885 1634 1648 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03529 1636 1635 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03528 1648 1639 1636 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03527 1885 1792 1641 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03526 1641 1868 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03525 1641 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03524 1626 1628 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03523 1628 1843 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03522 1885 1642 1628 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03521 1628 1836 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03520 1885 1850 1628 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03519 1629 1732 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03518 1885 1850 1631 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03517 1630 1631 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03516 1885 1642 1631 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03515 1631 1843 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03514 1732 1873 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03513 1885 1627 1732 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03512 1885 1736 1625 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03511 1757 1623 1625 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03510 1625 1624 1757 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03509 1885 1737 1622 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03508 1758 1622 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03507 1885 1736 1622 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03506 1622 1752 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03505 1885 1610 1615 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03504 1615 1614 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03503 1885 1613 1614 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03502 1621 1620 1737 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03501 1885 1619 1621 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03500 1751 1624 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03499 1885 1836 1612 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03498 1616 1612 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03497 1885 1611 1612 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03496 1612 1842 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03495 1605 1719 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03494 1885 1806 1606 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03493 1611 1605 1607 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03492 1607 1806 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03491 1607 1606 1611 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03490 1885 1719 1607 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03489 1712 1609 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03488 1609 1836 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03487 1885 1783 1609 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03486 1609 1806 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03485 1885 1719 1609 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03484 1885 1837 1608 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03483 1713 1608 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03482 1885 1783 1608 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03481 1608 1611 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03480 1885 1617 1702 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03479 1618 1732 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03478 1618 1615 1617 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03477 1617 1616 1618 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03476 1603 1601 1604 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03475 1885 1702 1603 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03474 1885 1599 1600 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03473 1600 1602 1601 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03472 1600 1806 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03471 1601 1842 1600 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03470 1885 1806 1602 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03469 1599 1842 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03468 1804 1598 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03467 1885 1595 1598 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03466 1653 1597 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03465 1885 1596 1597 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03464 1613 1806 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03463 1885 1873 1566 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03462 1567 1566 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03461 1885 1630 1566 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03460 1566 1875 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03459 1563 1562 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03458 1562 1873 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03457 1885 1630 1562 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03456 1562 1561 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03455 1885 1875 1562 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03454 1502 1792 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03453 1584 1587 1502 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03452 1589 1593 1584 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03451 1586 1593 1504 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03450 1504 1589 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03449 1505 1587 1586 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03448 1593 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03447 1885 1593 1587 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03446 1591 1592 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03445 1885 1591 1505 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03444 1885 1584 1792 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03443 1792 1584 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03442 1589 1586 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03441 1885 1641 1592 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03440 1501 1868 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03439 1592 1799 1501 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03438 1885 1629 1489 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03437 1559 1620 1489 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03436 1489 1557 1559 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03435 1490 1563 1557 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03434 1885 1845 1490 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03433 1486 1551 1549 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03432 1885 1703 1486 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03431 1553 1549 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03430 1548 1547 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03429 1547 1873 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03428 1885 1626 1547 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03427 1547 1561 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03426 1885 1875 1547 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03425 1574 1559 1488 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03424 1488 1840 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03423 1487 1845 1574 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03422 1885 1553 1487 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03421 1496 1620 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03420 1570 1576 1496 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03419 1575 1579 1570 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03418 1571 1579 1499 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03417 1499 1575 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03416 1498 1576 1571 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03415 1579 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03414 1885 1579 1576 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03413 1573 1574 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03412 1885 1573 1498 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03411 1885 1570 1620 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03410 1620 1570 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03409 1575 1571 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03408 1481 1868 1482 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03407 1885 1703 1481 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03406 1535 1548 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03405 1885 1540 1535 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03404 1480 1548 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03403 1885 1540 1480 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03402 1833 1542 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03401 1885 1551 1542 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03400 1542 1563 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03399 1540 1539 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03398 1885 1613 1539 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03397 1539 1719 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03396 1840 1703 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03395 1885 1534 1473 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03394 1472 1620 1474 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03393 1474 1736 1527 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03392 1473 1831 1472 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03391 1885 1845 1477 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03390 1477 1534 1476 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03389 1476 1533 1532 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03388 1624 1532 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03387 1475 1620 1533 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03386 1885 1535 1475 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03385 1524 1523 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03384 1885 1840 1523 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03383 1523 1527 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03382 1459 1806 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03381 1508 1511 1459 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03380 1510 1517 1508 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03379 1509 1517 1462 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03378 1462 1510 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03377 1461 1511 1509 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03376 1517 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03375 1885 1517 1511 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03374 1512 1513 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03373 1885 1512 1461 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03372 1885 1508 1806 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03371 1806 1508 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03370 1510 1509 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03369 1467 1833 1470 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03368 1885 1522 1467 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03367 1513 1518 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03366 1468 1470 1464 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03365 1468 1469 1885 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03364 1885 1703 1468 1885 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03363 1464 1604 1518 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03362 1518 1840 1468 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03361 1471 1613 1521 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03360 1885 1845 1471 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03359 1522 1521 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03358 1534 1752 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03357 1469 1522 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03356 1435 1433 1434 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03355 1885 1845 1435 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03354 1436 1434 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03353 1448 1447 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03352 1885 1868 1447 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03351 1447 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03350 1443 1436 1438 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03349 1438 1553 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03348 1437 1567 1443 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03347 1885 1436 1437 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03346 1449 1561 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03345 1450 1458 1449 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03344 1451 1457 1450 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03343 1453 1457 1452 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03342 1452 1451 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03341 1456 1458 1453 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03340 1457 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03339 1885 1457 1458 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03338 1455 1454 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03337 1885 1455 1456 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03336 1885 1450 1561 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03335 1561 1450 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03334 1451 1453 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03333 1418 1417 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03332 1420 1422 1418 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03331 1419 1427 1420 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03330 1425 1427 1424 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03329 1424 1419 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03328 1426 1422 1425 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03327 1427 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03326 1885 1427 1422 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03325 1423 1421 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03324 1885 1423 1426 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03323 1885 1420 1417 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03322 1417 1420 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03321 1419 1425 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03320 1885 1620 1428 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03319 1429 1433 1430 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03318 1430 1441 1627 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03317 1428 1779 1429 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03316 1885 1779 1440 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03315 1439 1561 1442 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03314 1442 1441 1444 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03313 1440 1840 1439 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03312 1431 1567 1432 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03311 1885 1845 1431 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03310 1885 1445 1454 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03309 1446 1443 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03308 1446 1444 1445 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03307 1445 1873 1446 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03306 1885 1540 1407 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03305 1407 1642 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03304 1407 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03303 1885 1845 1393 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03302 1396 1524 1395 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03301 1393 1411 1396 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03300 1885 1416 1415 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03299 1408 1415 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03298 1885 1410 1415 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03297 1415 1482 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03296 1885 1398 1421 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03295 1397 1395 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03294 1397 1405 1398 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03293 1398 1524 1397 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03292 1885 1411 1412 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03291 1414 1433 1413 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03290 1413 1736 1416 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03289 1412 1620 1414 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03288 1885 1480 1406 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03287 1406 1417 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03286 1406 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03285 1885 1875 1409 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03284 1410 1409 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03283 1885 1752 1409 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03282 1409 1842 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03281 1885 1406 1405 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03280 1404 1619 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03279 1405 1417 1404 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03278 1400 1736 1403 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03277 1401 1399 1400 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03276 1402 1417 1401 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03275 1885 1752 1402 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03274 1885 1403 1610 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03273 1885 1388 1390 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03272 1390 1389 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03271 1885 1448 1389 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03270 1885 1384 1387 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03269 1386 1385 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03268 1387 1390 1386 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03267 1394 1392 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03266 1885 1391 1392 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03265 1885 1385 1384 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03264 1384 1382 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03263 1384 1388 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03262 1373 1595 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03261 1374 1380 1373 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03260 1375 1381 1374 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03259 1378 1381 1377 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03258 1377 1375 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03257 1379 1380 1378 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03256 1381 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03255 1885 1381 1380 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03254 1376 1387 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03253 1885 1376 1379 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03252 1885 1374 1595 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03251 1595 1374 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03250 1375 1378 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03249 1885 1845 1388 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03248 1388 1383 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03247 1885 1595 1383 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03246 1353 1358 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03245 1885 1873 1358 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03244 1358 1875 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03243 1220 1385 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03242 1367 1315 1220 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03241 1369 1316 1367 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03240 1370 1316 1311 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03239 1311 1369 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03238 1310 1315 1370 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03237 1316 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03236 1885 1316 1315 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03235 1314 1313 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03234 1885 1314 1310 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03233 1885 1367 1385 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03232 1385 1367 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03231 1369 1370 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03230 1211 1873 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03229 1361 1304 1211 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03228 1363 1308 1361 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03227 1364 1308 1299 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03226 1299 1363 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03225 1302 1304 1364 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03224 1308 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03223 1885 1308 1304 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03222 1303 1448 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03221 1885 1303 1302 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03220 1885 1361 1873 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03219 1873 1361 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03218 1363 1364 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03217 1307 1306 1313 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03216 1885 1845 1307 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03215 1885 1853 1297 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03214 1297 1792 1296 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03213 1296 1298 1360 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03212 1441 1360 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03211 1885 1441 1290 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03210 1293 1703 1294 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03209 1294 1779 1295 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03208 1290 1868 1293 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03207 1298 1642 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03206 1289 1295 1359 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03205 1289 1432 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03204 1885 1703 1289 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03203 1359 1288 1289 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03202 1287 1359 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03201 1885 1354 1283 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03200 1283 1355 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03199 1283 1353 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03198 1551 1620 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03197 1885 1271 1341 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03196 1267 1341 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03195 1885 1268 1341 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03194 1341 1264 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03193 1885 1620 1280 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03192 1279 1613 1354 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03191 1280 1433 1279 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03190 1623 1281 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03189 1885 1283 1623 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03188 1277 1868 1350 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03187 1278 1433 1277 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03186 1276 1779 1278 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03185 1885 1274 1276 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03184 1885 1350 1619 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03183 1275 1407 1347 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03182 1272 1861 1275 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03181 1273 1792 1272 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03180 1885 1837 1273 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03179 1885 1347 1274 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03178 1885 1247 1329 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03177 1244 1329 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03176 1885 1240 1329 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03175 1329 1241 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03174 1885 1642 1250 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03173 1250 1385 1251 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03172 1251 1249 1330 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03171 1247 1330 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03170 1174 1391 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03169 1334 1262 1174 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03168 1335 1263 1334 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03167 1336 1263 1257 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03166 1257 1335 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03165 1256 1262 1336 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03164 1263 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03163 1885 1263 1262 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03162 1258 1267 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03161 1885 1258 1256 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03160 1885 1334 1391 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03159 1391 1334 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03158 1335 1336 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03157 1885 1845 1270 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03156 1270 1875 1269 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03155 1269 1385 1343 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03154 1271 1343 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03153 1261 1783 1338 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03152 1885 1391 1261 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03151 1268 1338 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03150 1248 1245 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03149 1885 1248 1246 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03148 1246 1783 1249 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03147 1153 1245 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03146 1319 1236 1153 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03145 1321 1239 1319 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03144 1322 1239 1231 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03143 1231 1321 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03142 1234 1236 1322 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03141 1239 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03140 1885 1239 1236 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03139 1235 1244 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03138 1885 1235 1234 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03137 1885 1319 1245 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03136 1245 1319 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03135 1321 1322 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03134 1885 1845 1254 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03133 1254 1837 1253 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03132 1253 1385 1333 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03131 1252 1333 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03130 1238 1783 1326 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03129 1885 1245 1238 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03128 1240 1326 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03127 1230 1318 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03126 1885 1245 1318 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03125 1214 1212 1215 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03124 1885 1213 1214 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03123 1885 1207 1210 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03122 1209 1208 1213 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03121 1210 1218 1209 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03120 1885 1215 1225 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03119 1225 1216 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03118 1225 1217 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03117 1219 1218 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03116 1224 1229 1219 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03115 1221 1227 1224 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03114 1223 1227 1222 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03113 1222 1221 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03112 1226 1229 1223 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03111 1227 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03110 1885 1227 1229 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03109 1228 1225 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03108 1885 1228 1226 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03107 1885 1224 1218 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03106 1218 1224 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03105 1221 1223 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03104 1885 1218 1206 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03103 1212 1206 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03102 1885 1783 1206 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03101 1206 1207 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03100 1355 1196 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03099 1196 1194 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03098 1885 1195 1196 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03097 1196 1626 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03096 1885 1411 1196 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03095 1199 1703 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03094 1198 1203 1199 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03093 1197 1205 1198 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03092 1202 1205 1204 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03091 1204 1197 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03090 1201 1203 1202 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03089 1205 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03088 1885 1205 1203 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03087 1200 1287 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03086 1885 1200 1201 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03085 1885 1198 1703 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03084 1703 1198 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03083 1197 1202 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03082 1433 1561 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03081 1411 1417 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03080 1288 1561 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03079 1885 1551 1288 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03078 1885 1191 1187 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03077 1192 1193 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03076 1192 1188 1191 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03075 1191 1408 1192 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03074 1195 1399 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03073 1885 1185 1188 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03072 1186 1274 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03071 1188 1399 1186 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03070 1885 1184 1185 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03069 1185 1399 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03068 1185 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03067 1184 1540 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03066 1885 1626 1184 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03065 1885 1845 1190 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03064 1189 1408 1193 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03063 1190 1195 1189 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03062 1885 1385 1157 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03061 1157 1154 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03060 1157 1155 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03059 1885 1155 1156 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03058 1156 1150 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03057 1156 1853 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03056 1885 1845 1155 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03055 1155 1152 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03054 1885 1596 1152 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03053 1173 1169 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03052 1172 1179 1173 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03051 1170 1182 1172 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03050 1178 1182 1171 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03049 1171 1170 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03048 1177 1179 1178 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03047 1182 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03046 1885 1182 1179 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03045 1176 1175 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03044 1885 1176 1177 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03043 1885 1172 1169 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03042 1169 1172 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03041 1170 1178 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03040 1158 1596 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03039 1159 1167 1158 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03038 1160 1165 1159 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03037 1162 1165 1163 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03036 1163 1160 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03035 1161 1167 1162 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03034 1165 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03033 1885 1165 1167 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03032 1166 1164 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03031 1885 1166 1161 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03030 1885 1159 1596 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03029 1596 1159 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03028 1160 1162 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03027 1151 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03026 1885 1831 1151 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03025 1180 1763 1183 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03024 1885 1845 1180 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03023 1181 1183 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03022 1507 1168 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03021 1885 1169 1168 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03020 1164 1157 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03019 1885 1156 1164 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03018 1148 1147 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03017 1885 1149 1147 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03016 1022 1101 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03015 1092 1100 1022 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03014 1093 1098 1092 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03013 1095 1098 1025 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03012 1025 1093 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03011 1024 1100 1095 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03010 1098 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03009 1885 1098 1100 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03008 1099 1097 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03007 1885 1099 1024 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03006 1885 1092 1101 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03005 1101 1092 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03004 1093 1095 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03003 1216 1109 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03002 1885 1105 1216 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03001 1885 1106 1109 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03000 1106 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02999 1885 1218 1032 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02998 1032 1104 1106 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02997 1885 1110 1038 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02996 1038 1112 1306 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02995 1038 1385 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02994 1306 1111 1038 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02993 1885 1385 1112 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02992 1110 1111 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02991 1028 1101 1102 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02990 1885 1104 1028 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02989 1103 1102 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02988 1885 1194 995 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02987 995 1385 998 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02986 998 1074 1076 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02985 1073 1076 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02984 1885 1433 1019 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02983 1019 1385 1018 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02982 1018 1089 1090 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02981 1088 1090 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02980 1014 1783 1089 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02979 1885 1087 1014 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02978 987 1783 1074 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02977 1885 1072 987 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02976 1002 1752 1281 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02975 1885 1845 1002 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02974 1194 1719 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02973 1069 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02972 1885 1068 1069 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02971 1001 1792 1077 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02970 1885 1845 1001 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02969 1075 1077 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02968 1005 1399 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02967 1080 1085 1005 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02966 1079 1086 1080 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02965 1084 1086 1009 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02964 1009 1079 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02963 1010 1085 1084 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02962 1086 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02961 1885 1086 1085 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02960 1081 1187 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02959 1885 1081 1010 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02958 1885 1080 1399 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02957 1399 1080 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02956 1079 1084 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02955 1885 1385 1065 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02954 1065 1069 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02953 1065 1067 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02952 1056 1057 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02951 1885 1087 1057 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02950 1175 1064 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02949 1885 1065 1175 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02948 1885 1075 1064 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02947 1064 1150 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02946 1064 1067 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02945 1885 1845 1067 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02944 1067 1060 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02943 1885 1169 1060 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02942 1885 1052 1054 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02941 1049 1054 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02940 1885 1051 1054 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02939 1054 1059 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02938 966 1783 1048 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02937 1885 1149 966 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02936 1051 1048 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02935 1885 1845 973 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02934 973 1703 976 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02933 976 1385 1055 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02932 1052 1055 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02931 958 1149 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02930 1040 1046 958 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02929 1041 1047 1040 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02928 1043 1047 961 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02927 961 1041 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02926 960 1046 1043 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02925 1047 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02924 1885 1047 1046 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02923 1042 1049 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02922 1885 1042 960 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02921 1885 1040 1149 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02920 1149 1040 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02919 1041 1043 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02918 1885 1031 1105 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02917 1105 1068 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02916 1885 1034 1105 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02915 1105 1035 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02914 1036 1037 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02913 1037 1033 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02912 1885 1034 1037 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02911 1037 1035 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02910 1885 1068 1037 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02909 1030 1036 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02908 1885 1029 1030 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02907 1885 1103 1027 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02906 1027 1030 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02905 1027 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02904 1885 1027 1097 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02903 1097 1023 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02902 1097 1026 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02901 1012 1011 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02900 1885 1029 1011 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02899 1011 1218 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02898 1016 1015 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02897 1885 1006 1007 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02896 1008 1007 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02895 1885 1012 1007 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02894 1007 1013 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02893 1026 1021 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02892 1885 1217 1021 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02891 1021 1020 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02890 1013 1017 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02889 1885 1068 1017 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02888 1017 1035 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02887 1006 1004 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02886 1885 1034 1004 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02885 1004 1015 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02884 1885 999 1000 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02883 1000 1088 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02882 1000 1003 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02881 989 1087 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02880 988 997 989 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02879 990 996 988 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02878 992 996 994 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02877 994 990 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02876 993 997 992 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02875 996 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02874 1885 996 997 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02873 991 1000 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02872 1885 991 993 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02871 1885 988 1087 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02870 1087 988 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02869 990 992 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02868 1885 1385 1059 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02867 1059 1034 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02866 1059 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02865 1003 1845 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02864 1885 1087 1003 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02863 979 931 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02862 1885 979 980 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02861 980 1783 982 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02860 986 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02859 1885 1551 986 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02858 1885 1806 983 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02857 983 1385 985 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02856 985 982 984 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02855 981 984 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02854 1885 1845 977 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02853 977 959 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02852 1885 962 959 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02851 975 974 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02850 1885 978 975 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02849 963 962 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02848 964 972 963 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02847 967 971 964 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02846 969 971 968 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02845 968 967 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02844 965 972 969 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02843 971 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02842 1885 971 972 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02841 970 975 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02840 1885 970 965 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02839 1885 964 962 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02838 962 964 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02837 967 969 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02836 1885 986 978 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02835 978 1150 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02834 978 977 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02833 957 956 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02832 1885 962 956 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02831 1885 1031 921 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02830 1033 921 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02829 1885 918 921 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02828 921 1218 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02827 1885 916 912 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02826 830 915 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02825 830 1036 916 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02824 916 914 830 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02823 1885 1783 915 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02822 823 1104 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02821 915 918 823 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02820 817 918 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02819 904 908 817 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02818 903 911 904 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02817 909 911 816 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02816 816 903 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02815 818 908 909 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02814 911 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02813 1885 911 908 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02812 907 906 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02811 1885 907 818 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02810 1885 904 918 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02809 918 904 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02808 903 909 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02807 1885 1217 906 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02806 906 898 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02805 1885 912 906 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02804 906 897 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02803 897 1207 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02802 1885 889 897 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02801 1885 1034 880 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02800 878 880 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02799 1885 1035 880 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02798 880 1068 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02797 1885 891 802 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02796 802 892 803 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02795 803 1016 893 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02794 894 893 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02793 1885 894 1020 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02792 1020 1101 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02791 1020 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02790 886 884 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02789 884 1034 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02788 1885 1031 884 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02787 884 1035 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02786 1885 1218 884 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02785 1885 874 872 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02784 872 1073 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02783 872 870 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02782 874 1385 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02781 1885 889 874 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02780 889 883 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02779 1885 918 883 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02778 883 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02777 999 1385 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02776 1885 879 999 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02775 1264 867 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02774 1885 1016 1264 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02773 1241 867 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02772 1885 891 1241 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02771 1885 1399 785 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02770 783 1385 857 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02769 785 1845 783 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02768 791 1072 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02767 863 866 791 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02766 860 869 863 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02765 862 869 794 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02764 794 860 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02763 797 866 862 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02762 869 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02761 1885 869 866 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02760 864 872 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02759 1885 864 797 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02758 1885 863 1072 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02757 1072 863 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02756 860 862 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02755 772 841 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02754 843 850 772 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02753 842 853 843 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02752 848 853 775 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02751 775 842 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02750 776 850 848 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02749 853 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02748 1885 853 850 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02747 846 845 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02746 1885 846 776 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02745 1885 843 841 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02744 841 843 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02743 842 848 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02742 856 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02741 1885 854 856 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02740 831 833 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02739 1885 841 833 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02738 1885 1151 839 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02737 839 1150 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02736 839 834 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02735 1885 1845 834 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02734 834 835 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02733 1885 841 835 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02732 1885 1385 974 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02731 974 856 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02730 974 977 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02729 845 838 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02728 1885 839 845 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02727 821 918 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02726 811 813 810 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02725 1885 812 811 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02724 1885 1101 819 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02723 820 821 825 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02722 825 822 824 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02721 819 828 820 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02720 1885 826 829 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02719 829 827 914 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02718 829 828 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02717 914 892 829 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02716 1885 828 827 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02715 826 892 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02714 1885 1035 1023 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02713 1023 815 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02712 1885 824 1023 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02711 1023 1068 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02710 756 757 800 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02709 1885 1207 756 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02708 805 800 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02707 804 892 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02706 1885 759 898 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02705 898 806 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02704 898 810 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02703 758 757 801 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02702 1885 894 758 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02701 822 801 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02700 814 813 815 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02699 1885 812 814 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02698 1885 918 807 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02697 809 804 808 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02696 808 805 806 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02695 807 1029 809 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02694 753 867 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02693 1885 1029 753 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02692 1034 812 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02691 751 867 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02690 1885 804 751 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02689 813 1218 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02688 1885 981 798 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02687 799 798 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02686 1885 796 798 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02685 798 751 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02684 870 1845 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02683 1885 1072 870 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02682 755 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02681 1885 813 755 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02680 784 931 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02679 788 782 784 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02678 789 786 788 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02677 787 786 790 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02676 790 789 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02675 792 782 787 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02674 786 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02673 1885 786 782 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02672 793 799 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02671 1885 793 792 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02670 1885 788 931 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02669 931 788 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02668 789 787 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02667 768 762 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02666 769 763 768 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02665 767 764 769 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02664 765 764 766 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02663 766 767 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02662 771 763 765 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02661 764 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02660 1885 764 763 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02659 770 781 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02658 1885 770 771 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02657 1885 769 762 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02656 762 769 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02655 767 765 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02654 746 1783 795 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02653 1885 931 746 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02652 796 795 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02651 1885 1752 779 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02650 778 1385 777 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02649 779 1845 778 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02648 1885 1252 780 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02647 781 780 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02646 1885 774 780 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02645 780 753 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02644 743 1783 773 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02643 1885 762 743 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02642 774 773 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02641 1885 1385 838 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02640 838 755 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02639 838 834 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02638 761 760 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02637 1885 931 760 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02636 642 1029 713 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02635 1885 716 642 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02634 711 713 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02633 719 918 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02632 1885 1029 719 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02631 1885 728 738 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02630 738 726 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02629 738 727 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02628 644 892 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02627 735 741 644 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02626 732 742 735 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02625 734 742 645 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02624 645 732 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02623 646 741 734 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02622 742 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02621 1885 742 741 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02620 740 738 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02619 1885 740 646 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02618 1885 735 892 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02617 892 735 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02616 732 734 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02615 1885 804 728 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02614 728 719 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02613 728 720 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02612 697 698 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02611 698 804 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02610 1885 1101 698 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02609 698 918 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02608 1885 710 698 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02607 643 804 717 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02606 1885 716 643 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02605 727 717 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02604 1885 709 716 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02603 641 707 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02602 641 886 709 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02601 709 1068 641 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02600 640 1104 706 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02599 1885 1845 640 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02598 707 706 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02597 1207 710 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02596 1885 1015 1207 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02595 1031 703 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02594 1885 1029 705 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02593 701 705 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02592 1885 1218 705 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02591 705 1015 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02590 691 692 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02589 1885 703 692 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02588 689 867 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02587 1885 689 638 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02586 638 1101 688 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02585 639 691 690 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02584 1885 695 639 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02583 1885 701 695 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02582 695 697 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02581 695 878 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02580 637 685 686 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02579 1885 707 637 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02578 687 686 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02577 631 673 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02576 667 675 631 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02575 666 674 667 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02574 671 674 633 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02573 633 666 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02572 632 675 671 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02571 674 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02570 1885 674 675 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02569 669 678 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02568 1885 669 632 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02567 1885 667 673 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02566 673 667 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02565 666 671 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02564 685 684 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02563 682 681 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02562 1885 685 681 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02561 681 867 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02560 1885 677 636 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02559 635 857 678 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02558 636 682 635 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02557 647 648 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02556 1885 762 648 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02555 628 1783 664 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02554 1885 661 628 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02553 626 661 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02552 653 658 626 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02551 655 662 653 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02550 652 662 625 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02549 625 655 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02548 627 658 652 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02547 662 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02546 1885 662 658 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02545 656 665 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02544 1885 656 627 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02543 1885 653 661 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02542 661 653 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02541 655 652 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02540 634 1783 677 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02539 1885 673 634 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02538 1885 688 629 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02537 630 777 665 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02536 629 664 630 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02535 1885 1029 623 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02534 623 624 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02533 1885 622 624 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02532 1885 711 617 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02531 617 616 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02530 617 623 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02529 1885 892 726 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02528 726 615 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02527 726 1207 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02526 614 1207 720 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02525 1885 619 614 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02524 621 618 620 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02523 1885 619 621 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02522 622 620 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02521 1885 604 605 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02520 607 892 606 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02519 605 891 607 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02518 1885 892 618 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02517 618 1015 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02516 618 710 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02515 612 1016 611 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02514 609 892 612 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02513 610 828 609 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02512 1885 813 610 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02511 1885 611 608 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02510 1885 828 616 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02509 616 615 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02508 616 618 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02507 879 613 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02506 1885 1035 613 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02505 613 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02504 594 684 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02503 595 603 594 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02502 597 602 595 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02501 600 602 599 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02500 599 597 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02499 598 603 600 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02498 602 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02497 1885 602 603 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02496 601 596 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02495 1885 601 598 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02494 1885 595 684 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02493 684 595 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02492 597 600 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02491 592 1101 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02490 1885 918 592 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02489 867 593 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02488 1885 1385 593 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02487 593 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02486 1885 583 585 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02485 587 684 586 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02484 586 588 589 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02483 585 584 587 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02482 1885 589 591 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02481 591 606 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02480 1885 1008 591 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02479 591 590 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02478 580 583 579 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02477 1885 684 580 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02476 576 560 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02475 1885 591 596 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02474 582 581 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02473 596 687 582 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02472 568 576 569 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02471 1885 1783 568 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02470 1885 1417 570 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02469 571 1385 572 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02468 570 569 571 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02467 574 575 573 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02466 1885 572 574 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02465 578 867 577 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02464 578 1845 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02463 1885 576 578 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02462 577 583 578 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02461 575 577 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02460 563 564 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02459 1885 567 563 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02458 1885 1385 564 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02457 564 566 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02456 564 565 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02455 1885 1181 567 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02454 567 1150 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02453 567 566 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02452 1150 1385 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02451 1885 1845 566 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02450 566 562 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02449 1885 561 562 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02448 537 1218 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02447 1885 1015 537 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02446 1208 541 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02445 1885 544 541 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02444 1029 828 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02443 459 544 545 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02442 1885 813 459 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02441 619 545 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02440 1885 534 458 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02439 457 537 535 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02438 458 533 457 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02437 460 828 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02436 554 557 460 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02435 553 558 554 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02434 552 558 461 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02433 461 553 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02432 462 557 552 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02431 558 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02430 1885 558 557 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02429 556 617 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02428 1885 556 462 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02427 1885 554 828 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02426 828 554 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02425 553 552 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02424 1885 526 524 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02423 524 527 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02422 1885 535 524 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02421 524 531 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02420 1885 604 452 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02419 454 892 453 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02418 453 891 531 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02417 452 828 454 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02416 1885 520 517 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02415 517 514 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02414 1885 532 517 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02413 517 513 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02412 1885 828 456 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02411 455 892 532 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02410 456 891 455 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02409 450 508 509 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02408 1885 517 450 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02407 1217 509 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02406 520 525 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02405 1885 1015 525 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02404 525 1218 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02403 451 534 513 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02402 1885 511 451 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02401 1885 1101 508 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02400 508 854 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02399 1885 501 508 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02398 508 918 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02397 1885 588 444 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02396 445 495 526 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02395 444 579 445 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02394 1885 524 500 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02393 448 690 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02392 500 498 448 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02391 449 592 590 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02390 1885 534 449 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02389 443 495 491 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02388 1885 1845 443 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02387 565 491 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02386 584 495 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02385 492 579 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02384 1885 492 442 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02383 442 565 501 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02382 1885 1845 447 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02381 447 1104 446 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02380 446 584 496 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02379 498 496 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02378 465 466 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02377 1885 1072 466 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02376 463 464 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02375 1885 673 464 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02374 439 495 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02373 482 490 439 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02372 484 488 482 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02371 485 488 441 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02370 441 484 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02369 440 490 485 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02368 488 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02367 1885 488 490 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02366 489 500 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02365 1885 489 440 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02364 1885 482 495 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02363 495 482 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02362 484 485 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02361 436 560 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02360 469 479 436 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02359 470 477 469 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02358 471 477 438 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02357 438 470 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02356 437 479 471 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02355 477 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02354 1885 477 479 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02353 478 573 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02352 1885 478 437 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02351 1885 469 560 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02350 560 469 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02349 470 471 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02348 403 419 514 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02347 1885 812 403 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02346 431 425 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02345 1885 424 431 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02344 426 1035 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02343 427 434 426 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02342 428 435 427 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02341 430 435 429 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02340 429 428 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02339 433 434 430 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02338 435 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02337 1885 435 434 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02336 432 431 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02335 1885 432 433 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02334 1885 427 1035 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02333 1035 427 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02332 428 430 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02331 1885 812 423 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02330 423 419 421 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02329 421 420 422 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02328 424 422 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02327 533 1101 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02326 1885 918 533 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02325 1885 396 414 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02324 394 402 396 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02323 395 608 394 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02322 398 391 395 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02321 398 397 1885 1885 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02320 1885 392 398 1885 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02319 398 400 1885 1885 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02318 396 393 398 1885 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_02317 401 407 400 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02316 1885 399 401 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02315 388 583 393 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02314 1885 1845 388 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02313 1885 812 404 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02312 404 511 406 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02311 406 419 405 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02310 402 405 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02309 420 418 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02308 392 695 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02307 1885 390 392 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02306 408 407 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02305 409 417 408 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02304 410 415 409 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02303 412 415 411 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02302 411 410 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02301 413 417 412 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02300 415 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02299 1885 415 417 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02298 416 414 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02297 1885 416 413 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02296 1885 409 407 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02295 407 409 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02294 410 412 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02293 583 407 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02292 1885 1101 391 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02291 391 918 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02290 1885 710 391 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02289 391 389 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02288 1885 854 703 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02287 703 390 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02286 703 381 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02285 389 384 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02284 384 390 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02283 1885 383 384 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02282 384 495 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02281 1885 854 384 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02280 387 583 386 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02279 1885 695 387 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02278 1885 377 378 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02277 377 390 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02276 1885 380 379 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02275 379 684 377 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02274 581 385 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02273 1885 386 385 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02272 385 389 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02271 383 382 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02270 1885 381 382 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02269 364 365 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02268 1885 661 365 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02267 1382 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02266 1885 374 1382 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02265 366 561 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02264 367 373 366 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02263 368 375 367 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02262 370 375 369 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02261 369 368 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02260 372 373 370 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02259 375 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02258 1885 375 373 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02257 371 563 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02256 1885 371 372 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02255 1885 367 561 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02254 561 367 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02253 368 370 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02252 1154 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02251 1885 376 1154 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02250 380 386 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02249 419 1035 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02248 1885 352 354 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02247 301 1104 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02246 354 1035 301 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02245 425 353 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02244 353 302 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02243 1885 1217 353 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02242 353 359 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02241 1885 354 353 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02240 307 306 358 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02239 1885 333 307 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02238 1885 812 359 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02237 359 419 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02236 359 358 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02235 302 306 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02234 1885 879 302 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02233 299 419 759 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02232 1885 511 299 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02231 296 345 347 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02230 297 812 296 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02229 298 511 297 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02228 1885 419 298 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02227 1885 347 544 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02226 891 710 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02225 1885 812 294 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02224 295 511 527 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02223 294 419 295 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02222 1885 604 291 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02221 291 534 293 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02220 293 292 344 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02219 345 344 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02218 757 346 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02217 1885 345 346 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02216 854 604 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02215 588 334 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02214 1885 292 334 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02213 1885 1845 290 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02212 289 534 418 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02211 290 854 289 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02210 327 324 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02209 1885 325 324 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02208 324 383 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02207 283 534 332 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02206 1885 588 283 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02205 333 332 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02204 1885 336 397 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02203 397 288 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02202 1885 534 288 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02201 1885 286 285 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02200 285 604 284 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02199 284 584 335 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02198 336 335 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02197 282 604 325 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02196 1885 495 282 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02195 1783 1845 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02194 1885 320 321 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02193 320 279 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02192 1885 327 280 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02191 280 534 320 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02190 276 278 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02189 1885 378 276 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02188 309 308 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02187 1885 561 308 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02186 196 534 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02185 310 273 196 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02184 315 274 310 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02183 313 274 270 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02182 270 315 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02181 269 273 313 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02180 274 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02179 1885 274 273 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02178 272 321 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02177 1885 272 269 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02176 1885 310 534 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02175 534 310 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02174 315 313 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02173 277 378 279 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02172 1885 1845 277 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02171 249 534 615 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02170 1885 1845 249 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02169 256 812 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02168 260 265 256 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02167 257 264 260 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02166 259 264 258 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02165 258 257 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02164 263 265 259 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02163 264 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02162 1885 264 265 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02161 262 261 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02160 1885 262 263 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02159 1885 260 812 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02158 812 260 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02157 257 259 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02156 1885 250 261 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02155 261 247 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02154 261 248 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02153 1885 253 255 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02152 255 254 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02151 1885 812 254 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02150 1885 812 250 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02149 250 615 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02148 250 306 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02147 267 891 266 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02146 1885 1845 267 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02145 248 244 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02144 1885 812 248 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02143 243 710 242 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02142 1885 399 243 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02141 252 251 352 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02140 1885 1845 252 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02139 1885 245 247 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02138 246 255 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02137 246 1035 245 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02136 245 854 246 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02135 241 240 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02134 240 812 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02133 1885 710 240 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02132 240 1035 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02131 1885 1015 240 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02130 1885 232 233 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02129 236 238 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02128 233 757 236 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02127 1885 235 234 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02126 239 233 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02125 239 418 235 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02124 235 238 239 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02123 1885 241 238 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02122 238 237 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02121 1885 511 237 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02120 232 244 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02119 1885 604 232 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02118 1885 1845 229 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02117 228 1104 244 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02116 229 383 228 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02115 231 286 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02114 1885 390 231 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02113 381 213 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02112 1885 211 213 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02111 213 376 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02110 188 190 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02109 1885 560 190 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02108 251 230 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02107 1885 390 230 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02106 230 383 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02105 1885 223 292 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02104 292 227 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02103 1885 226 227 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02102 216 604 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02101 217 225 216 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02100 218 224 217 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02099 221 224 220 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02098 220 218 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02097 222 225 221 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02096 224 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02095 1885 224 225 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02094 219 234 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02093 1885 219 222 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02092 1885 217 604 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02091 604 217 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02090 218 221 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02089 214 374 215 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02088 1885 226 214 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02087 286 215 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02086 1885 534 206 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02085 209 212 208 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02084 206 202 209 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02083 1885 276 203 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02082 203 200 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02081 203 1783 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02080 210 325 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02079 1885 210 207 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02078 207 226 212 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02077 205 208 204 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02076 1885 203 205 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02075 191 189 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02074 192 198 191 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02073 193 201 192 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02072 195 201 194 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02071 194 193 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02070 199 198 195 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02069 201 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02068 1885 201 198 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02067 197 204 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02066 1885 197 199 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02065 1885 192 189 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02064 189 192 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02063 193 195 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02062 157 266 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02061 1885 155 157 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02060 1885 157 150 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02059 150 148 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02058 150 1217 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02057 1885 1015 155 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02056 155 1068 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02055 155 251 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02054 152 306 253 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02053 1885 333 152 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02052 123 534 124 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02051 1885 122 123 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02050 125 124 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02049 1885 137 144 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02048 61 134 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02047 61 135 137 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02046 137 1015 61 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02045 128 1068 130 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02044 1885 1845 128 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02043 56 131 132 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02042 56 352 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02041 1885 1068 56 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02040 132 130 56 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02039 135 132 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02038 1885 231 148 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02037 148 125 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02036 148 242 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02035 65 1015 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02034 139 146 65 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02033 140 147 139 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02032 143 147 68 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02031 68 140 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02030 67 146 143 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02029 147 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02028 1885 147 146 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02027 145 144 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02026 1885 145 67 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02025 1885 139 1015 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02024 1015 139 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02023 140 143 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02022 118 111 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02021 1885 390 111 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02020 111 1068 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02019 1885 399 119 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02018 119 118 120 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02017 120 1015 121 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02016 117 121 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02015 112 109 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02014 1885 226 109 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02013 109 278 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02012 131 112 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02011 1885 390 131 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02010 1885 1217 134 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02009 115 114 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02008 134 117 115 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02007 211 96 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02006 102 376 101 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02005 101 104 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02004 100 333 102 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02003 1885 122 100 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02002 390 534 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02001 96 189 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02000 1885 93 96 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01999 278 97 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01998 1885 211 97 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01997 19 226 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01996 85 92 19 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01995 86 90 85 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01994 89 90 23 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01993 23 86 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01992 22 92 89 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01991 90 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01990 1885 90 92 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01989 91 102 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01988 1885 91 22 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01987 1885 85 226 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01986 226 85 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01985 86 89 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01984 1885 1845 106 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01983 106 278 105 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01982 105 1104 107 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01981 104 107 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01980 202 94 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01979 1885 96 94 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01978 1885 534 98 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01977 114 226 98 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01976 98 189 114 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01975 374 189 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01974 1885 79 82 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01973 82 81 83 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01972 82 80 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01971 83 187 82 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01970 1885 80 81 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01969 79 187 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01968 306 122 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01967 1885 710 306 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01966 122 52 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01965 1885 1068 52 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01964 52 1015 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01963 66 710 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01962 73 75 66 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01961 69 76 73 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01960 71 76 70 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01959 70 69 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01958 72 75 71 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01957 76 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01956 1885 76 75 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01955 74 150 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01954 1885 74 72 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01953 1885 73 710 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01952 710 73 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01951 69 71 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01950 78 83 77 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01949 1885 1845 78 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01948 1068 511 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01947 54 53 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01946 55 64 54 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01945 57 62 55 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01944 59 62 60 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01943 60 57 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01942 58 64 59 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01941 62 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01940 1885 62 64 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01939 63 77 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01938 1885 63 58 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01937 1885 55 53 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01936 53 55 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01935 57 59 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01934 42 511 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01933 43 51 42 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01932 44 50 43 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01931 45 50 47 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01930 47 44 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01929 46 51 45 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01928 50 1881 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01927 1885 50 51 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01926 49 48 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01925 1885 49 46 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01924 1885 43 511 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01923 511 43 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01922 44 45 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01921 1885 41 48 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01920 40 38 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01919 40 511 41 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01918 41 39 40 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01917 1104 32 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01916 1885 534 32 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01915 32 80 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01914 1885 34 37 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01913 38 37 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01912 1885 118 37 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01911 37 226 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01910 1885 1845 36 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01909 35 1104 39 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01908 36 112 35 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01907 34 33 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01906 1885 223 33 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01905 1885 53 27 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01904 1885 27 93 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01903 93 27 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01902 1885 27 93 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01901 93 27 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01900 399 31 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01899 1885 30 31 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01898 80 28 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01897 1885 93 28 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01896 1885 53 24 1885 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_01895 24 53 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01894 376 226 1885 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01893 200 374 1885 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01892 1885 26 200 1885 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01891 29 30 223 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01890 1885 374 29 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01889 26 25 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01888 1885 24 25 1885 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01887 20 24 21 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01886 1885 1845 20 1885 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01885 30 21 1885 1885 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01884 1777 1871 1863 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01883 1803 1861 1777 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01882 1863 1872 1864 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01881 1803 1864 1781 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01880 1781 1872 1867 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01879 1867 1871 1782 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01878 1872 1871 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01877 1803 1881 1871 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01876 1782 1870 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01875 1803 1869 1870 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01874 1861 1863 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01873 1803 1863 1861 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01872 1864 1867 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01871 1791 1886 1876 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01870 1803 1875 1791 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01869 1876 1884 1877 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01868 1803 1877 1796 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01867 1796 1884 1879 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01866 1879 1886 1802 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01865 1884 1886 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01864 1803 1881 1886 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01863 1802 1883 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01862 1803 1880 1883 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01861 1875 1876 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01860 1803 1876 1875 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01859 1877 1879 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01858 1803 1856 1769 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01857 1769 1873 1855 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01856 1858 1847 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01855 1847 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01854 1803 1843 1847 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01853 1857 1854 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01852 1854 1853 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01851 1803 1856 1854 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01850 1803 1873 1775 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01849 1775 1858 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01848 1869 1868 1775 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01847 1775 1857 1869 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01846 1851 1875 1762 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01845 1803 1851 1856 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01844 1762 1850 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01843 1803 1873 1868 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01842 1849 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01841 1803 1846 1849 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01840 1853 1839 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01839 1839 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01838 1803 1861 1839 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01837 1832 1835 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01836 1835 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01835 1803 1833 1835 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01834 1803 1837 1836 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01833 1803 1861 1843 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01832 1808 1806 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01831 1803 1837 1805 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01830 1686 1805 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01829 1809 1808 1686 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01828 1692 1837 1809 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01827 1803 1806 1692 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01826 1803 1833 1711 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01825 1711 1840 1818 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01824 1803 1842 1831 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01823 1841 1842 1747 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01822 1803 1841 1846 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01821 1747 1840 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01820 1810 1809 1695 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01819 1803 1810 1813 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01818 1695 1842 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01817 1721 1829 1822 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01816 1803 1837 1721 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01815 1822 1830 1823 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01814 1803 1823 1727 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01813 1727 1830 1828 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01812 1828 1829 1726 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01811 1830 1829 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01810 1803 1881 1829 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01809 1726 1826 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01808 1803 1824 1826 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01807 1837 1822 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01806 1803 1822 1837 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01805 1823 1828 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01804 1820 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01803 1803 1836 1820 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01802 1803 1815 1824 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01801 1803 1813 1706 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01800 1706 1812 1803 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01799 1815 1820 1710 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01798 1710 1818 1803 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01797 1706 1814 1815 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01796 1811 1837 1701 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01795 1803 1811 1812 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01794 1701 1831 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01793 1803 1792 1850 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01792 1798 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01791 1800 1797 1799 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01790 1803 1798 1800 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01789 1801 1861 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01788 1803 1792 1794 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01787 1795 1794 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01786 1797 1801 1795 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01785 1793 1792 1797 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01784 1803 1861 1793 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01783 1880 1790 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01782 1803 1787 1790 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01781 1789 1788 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01780 1790 1873 1789 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01779 1756 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01778 1803 1846 1756 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01777 1780 1779 1788 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01776 1788 1799 1780 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01775 1780 1778 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01774 1803 1875 1779 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01773 1803 1786 1787 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01772 1784 1868 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01771 1785 1875 1784 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01770 1786 1783 1785 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01769 1776 1850 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01768 1776 1858 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01767 1803 1875 1776 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01766 1803 1776 1778 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01765 1803 1763 1736 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01764 1803 1760 1770 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01763 1803 1757 1761 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01762 1761 1758 1803 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01761 1760 1849 1759 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01760 1759 1763 1803 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01759 1761 1846 1760 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01758 1803 1753 1749 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01757 1803 1750 1754 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01756 1754 1751 1803 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01755 1753 1756 1755 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01754 1755 1752 1803 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01753 1754 1846 1753 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01752 1764 1774 1768 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01751 1803 1763 1764 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01750 1768 1773 1765 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01749 1803 1765 1766 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01748 1766 1773 1767 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01747 1767 1774 1771 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01746 1773 1774 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01745 1803 1881 1774 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01744 1771 1772 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01743 1803 1770 1772 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01742 1763 1768 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01741 1803 1768 1763 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01740 1765 1767 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01739 1803 1737 1738 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01738 1750 1738 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01737 1803 1752 1750 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01736 1714 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01735 1803 1715 1714 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01734 1803 1732 1735 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01733 1735 1842 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01732 1733 1831 1735 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01731 1735 1832 1733 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01730 1803 1707 1715 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01729 1708 1840 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01728 1709 1842 1708 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01727 1707 1833 1709 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01726 1720 1734 1725 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01725 1803 1719 1720 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01724 1725 1730 1722 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01723 1803 1722 1723 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01722 1723 1730 1724 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01721 1724 1734 1731 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01720 1730 1734 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01719 1803 1881 1734 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01718 1731 1729 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01717 1803 1728 1729 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01716 1719 1725 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01715 1803 1725 1719 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01714 1722 1724 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01713 1803 1716 1728 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01712 1803 1712 1717 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01711 1717 1713 1803 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01710 1716 1714 1718 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01709 1718 1719 1803 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01708 1717 1715 1716 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01707 1700 1705 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01706 1803 1696 1705 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01705 1704 1733 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01704 1705 1840 1704 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01703 1814 1702 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01702 1803 1703 1814 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01701 1739 1748 1742 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01700 1803 1752 1739 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01699 1742 1743 1740 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01698 1803 1740 1741 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01697 1741 1743 1745 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01696 1745 1748 1746 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01695 1743 1748 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01694 1803 1881 1748 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01693 1746 1744 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01692 1803 1749 1744 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01691 1752 1742 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01690 1803 1742 1752 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01689 1740 1745 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01688 1803 1699 1696 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01687 1697 1703 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01686 1698 1842 1697 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01685 1699 1783 1698 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01684 1684 1694 1685 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01683 1803 1842 1684 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01682 1685 1693 1687 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01681 1803 1687 1689 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01680 1689 1693 1690 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01679 1690 1694 1691 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01678 1693 1694 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01677 1803 1881 1694 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01676 1691 1688 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01675 1803 1700 1688 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01674 1842 1685 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01673 1803 1685 1842 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01672 1687 1690 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01671 1803 1783 1569 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01670 1569 1855 1568 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01669 1568 1642 1634 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01668 1640 1861 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01667 1803 1642 1637 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01666 1578 1637 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01665 1639 1640 1578 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01664 1580 1642 1639 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01663 1803 1861 1580 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01662 1585 1652 1644 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01661 1803 1642 1585 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01660 1644 1651 1645 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01659 1803 1645 1590 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01658 1590 1651 1646 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01657 1646 1652 1594 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01656 1651 1652 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01655 1803 1881 1652 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01654 1594 1649 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01653 1803 1648 1649 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01652 1642 1644 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01651 1803 1644 1642 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01650 1645 1646 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01649 1635 1633 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01648 1633 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01647 1803 1855 1633 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01646 1572 1635 1648 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01645 1648 1639 1572 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01644 1572 1634 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01643 1803 1783 1583 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01642 1583 1792 1582 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01641 1582 1868 1641 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01640 1555 1836 1552 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01639 1803 1843 1556 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01638 1552 1850 1628 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01637 1556 1642 1555 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01636 1803 1628 1626 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01635 1803 1732 1629 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01634 1803 1631 1630 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01633 1564 1850 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01632 1565 1843 1564 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01631 1631 1642 1565 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01630 1803 1873 1560 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01629 1560 1627 1732 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01628 1803 1623 1550 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01627 1550 1624 1757 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01626 1757 1736 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01625 1803 1622 1758 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01624 1545 1737 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01623 1546 1752 1545 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01622 1622 1736 1546 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01621 1614 1613 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01620 1538 1610 1615 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01619 1803 1614 1538 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01618 1737 1619 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01617 1803 1620 1737 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01616 1803 1624 1751 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01615 1803 1612 1616 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01614 1536 1836 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01613 1537 1842 1536 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01612 1612 1611 1537 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01611 1606 1806 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01610 1803 1719 1605 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01609 1519 1605 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01608 1611 1606 1519 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01607 1520 1719 1611 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01606 1803 1806 1520 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01605 1530 1806 1529 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01604 1803 1836 1531 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01603 1529 1719 1609 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01602 1531 1783 1530 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01601 1803 1609 1712 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01600 1803 1608 1713 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01599 1525 1837 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01598 1526 1611 1525 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01597 1608 1783 1526 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01596 1702 1617 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01595 1803 1732 1617 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01594 1541 1615 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01593 1617 1616 1541 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01592 1604 1702 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01591 1803 1601 1604 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01590 1803 1806 1516 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01589 1516 1599 1601 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01588 1601 1602 1515 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01587 1515 1842 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01586 1803 1842 1599 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01585 1602 1806 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01584 1803 1598 1804 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01583 1598 1595 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01582 1803 1597 1653 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01581 1597 1596 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01580 1803 1806 1613 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01579 1803 1566 1567 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01578 1495 1873 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01577 1494 1875 1495 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01576 1566 1630 1494 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01575 1492 1561 1491 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01574 1803 1873 1493 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01573 1491 1875 1562 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01572 1493 1630 1492 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01571 1803 1562 1563 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01570 1503 1593 1584 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01569 1803 1792 1503 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01568 1584 1587 1589 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01567 1803 1589 1588 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01566 1588 1587 1586 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01565 1586 1593 1506 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01564 1587 1593 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01563 1803 1881 1593 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01562 1506 1591 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01561 1803 1592 1591 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01560 1792 1584 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01559 1803 1584 1792 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01558 1589 1586 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01557 1581 1868 1592 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01556 1592 1799 1581 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01555 1581 1641 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01554 1803 1620 1558 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01553 1558 1557 1559 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01552 1559 1629 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01551 1557 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01550 1803 1563 1557 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01549 1553 1549 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01548 1549 1703 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01547 1803 1551 1549 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01546 1483 1561 1484 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01545 1803 1873 1485 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01544 1484 1875 1547 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01543 1485 1626 1483 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01542 1803 1547 1548 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01541 1803 1553 1554 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01540 1554 1845 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01539 1574 1559 1554 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01538 1554 1840 1574 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01537 1497 1579 1570 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01536 1803 1620 1497 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01535 1570 1576 1575 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01534 1803 1575 1577 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01533 1577 1576 1571 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01532 1571 1579 1500 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01531 1576 1579 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01530 1803 1881 1579 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01529 1500 1573 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01528 1803 1574 1573 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01527 1620 1570 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01526 1803 1570 1620 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01525 1575 1571 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01524 1482 1703 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01523 1803 1868 1482 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01522 1803 1548 1478 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01521 1478 1540 1535 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01520 1803 1548 1479 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01519 1479 1540 1480 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01518 1542 1563 1544 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01517 1803 1542 1833 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01516 1544 1551 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01515 1539 1719 1543 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01514 1803 1539 1540 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01513 1543 1613 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01512 1803 1703 1840 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01511 1527 1534 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01510 1803 1736 1527 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01509 1803 1831 1527 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01508 1527 1620 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01507 1532 1533 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01506 1532 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01505 1803 1534 1532 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01504 1803 1532 1624 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01503 1533 1535 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01502 1803 1620 1533 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01501 1523 1527 1528 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01500 1803 1523 1524 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01499 1528 1840 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01498 1460 1517 1508 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01497 1803 1806 1460 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01496 1508 1511 1510 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01495 1803 1510 1514 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01494 1514 1511 1509 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01493 1509 1517 1463 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01492 1511 1517 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01491 1803 1881 1517 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01490 1463 1512 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01489 1803 1513 1512 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01488 1806 1508 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01487 1803 1508 1806 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01486 1510 1509 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01485 1470 1522 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01484 1803 1833 1470 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01483 1803 1518 1513 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01482 1803 1604 1466 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01481 1466 1470 1803 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01480 1518 1469 1465 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01479 1465 1703 1803 1803 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01478 1466 1840 1518 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01477 1522 1521 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01476 1521 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01475 1803 1613 1521 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01474 1803 1752 1534 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01473 1803 1522 1469 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01472 1436 1434 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01471 1434 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01470 1803 1433 1434 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01469 1447 1783 1366 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01468 1803 1447 1448 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01467 1366 1868 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01466 1803 1436 1362 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01465 1362 1567 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01464 1443 1436 1362 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01463 1362 1553 1443 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01462 1368 1457 1450 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01461 1803 1561 1368 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01460 1450 1458 1451 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01459 1803 1451 1371 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01458 1371 1458 1453 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01457 1453 1457 1372 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01456 1458 1457 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01455 1803 1881 1457 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01454 1372 1455 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01453 1803 1454 1455 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01452 1561 1450 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01451 1803 1450 1561 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01450 1451 1453 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01449 1352 1427 1420 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01448 1803 1417 1352 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01447 1420 1422 1419 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01446 1803 1419 1356 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01445 1356 1422 1425 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01444 1425 1427 1357 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01443 1422 1427 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01442 1803 1881 1427 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01441 1357 1423 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01440 1803 1421 1423 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01439 1417 1420 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01438 1803 1420 1417 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01437 1419 1425 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01436 1627 1620 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01435 1803 1441 1627 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01434 1803 1779 1627 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01433 1627 1433 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01432 1444 1779 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01431 1803 1441 1444 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01430 1803 1840 1444 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01429 1444 1561 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01428 1432 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01427 1803 1567 1432 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01426 1454 1445 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01425 1803 1443 1445 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01424 1365 1444 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01423 1445 1873 1365 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01422 1803 1783 1346 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01421 1346 1540 1345 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01420 1345 1642 1407 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01419 1803 1411 1395 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01418 1395 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01417 1395 1524 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01416 1803 1415 1408 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01415 1349 1416 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01414 1351 1482 1349 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01413 1415 1410 1351 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01412 1421 1398 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01411 1803 1395 1398 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01410 1337 1405 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01409 1398 1524 1337 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01408 1416 1411 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01407 1803 1736 1416 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01406 1803 1620 1416 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01405 1416 1433 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01404 1803 1783 1342 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01403 1342 1480 1340 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01402 1340 1417 1406 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01401 1803 1409 1410 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01400 1344 1875 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01399 1348 1842 1344 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01398 1409 1752 1348 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01397 1339 1619 1405 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01396 1405 1417 1339 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01395 1339 1406 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01394 1403 1752 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01393 1803 1736 1403 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01392 1803 1417 1403 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01391 1403 1399 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01390 1610 1403 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01389 1389 1448 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01388 1332 1388 1390 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01387 1803 1389 1332 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01386 1331 1385 1387 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01385 1387 1390 1331 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01384 1331 1384 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01383 1803 1392 1394 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01382 1392 1391 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01381 1803 1388 1328 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01380 1328 1385 1327 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01379 1327 1382 1384 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01378 1320 1381 1374 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01377 1803 1595 1320 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01376 1374 1380 1375 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01375 1803 1375 1324 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01374 1324 1380 1378 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01373 1378 1381 1323 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01372 1380 1381 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01371 1803 1881 1381 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01370 1323 1376 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01369 1803 1387 1376 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01368 1595 1374 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01367 1803 1374 1595 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01366 1375 1378 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01365 1383 1595 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01364 1325 1845 1388 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01363 1803 1383 1325 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01362 1358 1875 1286 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01361 1803 1358 1353 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01360 1286 1873 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01359 1309 1316 1367 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01358 1803 1385 1309 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01357 1367 1315 1369 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01356 1803 1369 1312 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01355 1312 1315 1370 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01354 1370 1316 1317 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01353 1315 1316 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01352 1803 1881 1316 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01351 1317 1314 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01350 1803 1313 1314 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01349 1385 1367 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01348 1803 1367 1385 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01347 1369 1370 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01346 1300 1308 1361 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01345 1803 1873 1300 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01344 1361 1304 1363 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01343 1803 1363 1301 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01342 1301 1304 1364 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01341 1364 1308 1305 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01340 1304 1308 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01339 1803 1881 1308 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01338 1305 1303 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01337 1803 1448 1303 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01336 1873 1361 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01335 1803 1361 1873 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01334 1363 1364 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01333 1313 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01332 1803 1306 1313 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01331 1360 1298 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01330 1360 1853 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01329 1803 1792 1360 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01328 1803 1360 1441 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01327 1295 1441 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01326 1803 1779 1295 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01325 1803 1868 1295 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01324 1295 1703 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01323 1803 1642 1298 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01322 1292 1295 1359 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01321 1803 1288 1292 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01320 1291 1432 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01319 1359 1703 1291 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01318 1803 1359 1287 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01317 1803 1353 1284 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01316 1284 1354 1285 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01315 1285 1355 1283 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01314 1803 1620 1551 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01313 1803 1341 1267 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01312 1265 1271 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01311 1266 1264 1265 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01310 1341 1268 1266 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01309 1803 1433 1354 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01308 1354 1620 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01307 1354 1613 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01306 1803 1281 1282 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01305 1282 1283 1623 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01304 1350 1274 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01303 1803 1868 1350 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01302 1803 1779 1350 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01301 1350 1433 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01300 1619 1350 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01299 1347 1837 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01298 1803 1407 1347 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01297 1803 1792 1347 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01296 1347 1861 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01295 1274 1347 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01294 1803 1329 1244 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01293 1242 1247 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01292 1243 1241 1242 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01291 1329 1240 1243 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01290 1330 1249 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01289 1330 1642 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01288 1803 1385 1330 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01287 1803 1330 1247 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01286 1255 1263 1334 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01285 1803 1391 1255 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01284 1334 1262 1335 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01283 1803 1335 1259 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01282 1259 1262 1336 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01281 1336 1263 1260 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01280 1262 1263 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01279 1803 1881 1263 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01278 1260 1258 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01277 1803 1267 1258 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01276 1391 1334 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01275 1803 1334 1391 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01274 1335 1336 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01273 1343 1385 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01272 1343 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01271 1803 1875 1343 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01270 1803 1343 1271 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01269 1268 1338 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01268 1338 1391 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01267 1803 1783 1338 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01266 1803 1245 1248 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01265 1249 1248 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01264 1803 1783 1249 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01263 1232 1239 1319 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01262 1803 1245 1232 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01261 1319 1236 1321 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01260 1803 1321 1233 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01259 1233 1236 1322 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01258 1322 1239 1237 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01257 1236 1239 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01256 1803 1881 1239 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01255 1237 1235 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01254 1803 1244 1235 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01253 1245 1319 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01252 1803 1319 1245 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01251 1321 1322 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01250 1333 1385 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01249 1333 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01248 1803 1837 1333 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01247 1803 1333 1252 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01246 1240 1326 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01245 1326 1245 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01244 1803 1783 1326 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01243 1803 1318 1230 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01242 1318 1245 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01241 1215 1213 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01240 1803 1212 1215 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01239 1803 1218 1213 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01238 1213 1207 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01237 1213 1208 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01236 1803 1217 1143 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01235 1143 1215 1142 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01234 1142 1216 1225 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01233 1144 1227 1224 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01232 1803 1218 1144 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01231 1224 1229 1221 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01230 1803 1221 1145 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01229 1145 1229 1223 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01228 1223 1227 1146 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01227 1229 1227 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01226 1803 1881 1227 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01225 1146 1228 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01224 1803 1225 1228 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01223 1218 1224 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01222 1803 1224 1218 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01221 1221 1223 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01220 1803 1206 1212 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01219 1141 1218 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01218 1140 1207 1141 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01217 1206 1783 1140 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01216 1135 1626 1134 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01215 1803 1194 1133 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01214 1134 1411 1196 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01213 1133 1195 1135 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01212 1803 1196 1355 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01211 1137 1205 1198 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01210 1803 1703 1137 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01209 1198 1203 1197 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01208 1803 1197 1138 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01207 1138 1203 1202 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01206 1202 1205 1139 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01205 1203 1205 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01204 1803 1881 1205 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01203 1139 1200 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01202 1803 1287 1200 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01201 1703 1198 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01200 1803 1198 1703 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01199 1197 1202 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01198 1803 1561 1433 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01197 1803 1417 1411 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01196 1803 1561 1136 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01195 1136 1551 1288 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01194 1187 1191 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01193 1803 1193 1191 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01192 1132 1188 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01191 1191 1408 1132 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01190 1803 1399 1195 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01189 1131 1274 1188 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01188 1188 1399 1131 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01187 1131 1185 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01186 1803 1783 1130 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01185 1130 1184 1129 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01184 1129 1399 1185 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01183 1803 1540 1128 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01182 1128 1626 1184 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01181 1803 1195 1193 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01180 1193 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01179 1193 1408 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01178 1803 1155 1120 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01177 1120 1385 1119 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01176 1119 1154 1157 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01175 1803 1853 1118 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01174 1118 1155 1117 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01173 1117 1150 1156 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01172 1152 1596 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01171 1115 1845 1155 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01170 1803 1152 1115 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01169 1126 1182 1172 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01168 1803 1169 1126 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01167 1172 1179 1170 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01166 1803 1170 1125 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01165 1125 1179 1178 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01164 1178 1182 1127 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01163 1179 1182 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01162 1803 1881 1182 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01161 1127 1176 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01160 1803 1175 1176 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01159 1169 1172 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01158 1803 1172 1169 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01157 1170 1178 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01156 1122 1165 1159 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01155 1803 1596 1122 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01154 1159 1167 1160 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01153 1803 1160 1123 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01152 1123 1167 1162 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01151 1162 1165 1124 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01150 1167 1165 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01149 1803 1881 1165 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01148 1124 1166 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01147 1803 1164 1166 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01146 1596 1159 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01145 1803 1159 1596 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01144 1160 1162 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01143 1803 1783 1116 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01142 1116 1831 1151 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01141 1181 1183 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01140 1183 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01139 1803 1763 1183 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01138 1803 1168 1507 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01137 1168 1169 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01136 1803 1157 1121 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01135 1121 1156 1164 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01134 1803 1147 1148 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01133 1147 1149 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01132 1091 1098 1092 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01131 1803 1101 1091 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01130 1092 1100 1093 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01129 1803 1093 1094 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01128 1094 1100 1095 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01127 1095 1098 1096 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01126 1100 1098 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01125 1803 1881 1098 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01124 1096 1099 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01123 1803 1097 1099 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01122 1101 1092 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01121 1803 1092 1101 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01120 1093 1095 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01119 1803 1109 1107 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01118 1107 1105 1216 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01117 1106 1218 1108 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01116 1108 1104 1106 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01115 1803 1783 1108 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01114 1109 1106 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01113 1803 1385 1114 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01112 1114 1110 1306 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01111 1306 1112 1113 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01110 1113 1111 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01109 1803 1111 1110 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01108 1112 1385 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01107 1103 1102 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01106 1102 1104 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01105 1803 1101 1102 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01104 1076 1074 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01103 1076 1194 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01102 1803 1385 1076 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01101 1803 1076 1073 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01100 1090 1089 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01099 1090 1433 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01098 1803 1385 1090 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01097 1803 1090 1088 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01096 1089 1087 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01095 1803 1783 1089 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01094 1074 1072 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01093 1803 1783 1074 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01092 1281 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01091 1803 1752 1281 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01090 1803 1719 1194 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01089 1803 1783 1071 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01088 1071 1068 1069 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01087 1075 1077 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01086 1077 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01085 1803 1792 1077 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01084 1078 1086 1080 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01083 1803 1399 1078 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01082 1080 1085 1079 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01081 1803 1079 1082 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01080 1082 1085 1084 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01079 1084 1086 1083 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01078 1085 1086 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01077 1803 1881 1086 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01076 1083 1081 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01075 1803 1187 1081 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01074 1399 1080 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01073 1803 1080 1399 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01072 1079 1084 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01071 1803 1067 1070 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01070 1070 1385 1066 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01069 1066 1069 1065 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01068 1803 1057 1056 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01067 1057 1087 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01066 1803 1064 1063 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01065 1063 1065 1175 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01064 1803 1067 1062 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01063 1062 1075 1061 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01062 1061 1150 1064 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01061 1060 1169 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01060 1058 1845 1067 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01059 1803 1060 1058 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01058 1803 1054 1049 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01057 1050 1052 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01056 1053 1059 1050 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01055 1054 1051 1053 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01054 1051 1048 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01053 1048 1149 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01052 1803 1783 1048 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01051 1055 1385 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01050 1055 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01049 1803 1703 1055 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01048 1803 1055 1052 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01047 1039 1047 1040 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01046 1803 1149 1039 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01045 1040 1046 1041 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01044 1803 1041 1044 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01043 1044 1046 1043 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01042 1043 1047 1045 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01041 1046 1047 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01040 1803 1881 1047 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01039 1045 1042 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01038 1803 1049 1042 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01037 1149 1040 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01036 1803 1040 1149 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01035 1041 1043 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01034 1803 1035 952 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01033 952 1031 951 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01032 951 1068 950 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01031 950 1034 1105 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01030 953 1035 955 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01029 1803 1033 954 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01028 955 1068 1037 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01027 954 1034 953 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01026 1803 1037 1036 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01025 1803 1036 949 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01024 949 1029 1030 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01023 1803 1783 947 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01022 947 1103 948 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01021 948 1030 1027 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01020 1803 1026 946 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01019 946 1027 945 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01018 945 1023 1097 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01017 1011 1218 942 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01016 1803 1011 1012 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01015 942 1029 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01014 1803 1015 1016 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01013 1803 1007 1008 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01012 940 1006 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01011 941 1013 940 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01010 1007 1012 941 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01009 1021 1020 944 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01008 1803 1021 1026 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01007 944 1217 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01006 1017 1035 943 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01005 1803 1017 1013 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01004 943 1068 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01003 1004 1015 939 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01002 1803 1004 1006 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01001 939 1034 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01000 1803 1003 937 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00999 937 999 936 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00998 936 1088 1000 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00997 933 996 988 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00996 1803 1087 933 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00995 988 997 990 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00994 1803 990 934 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00993 934 997 992 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00992 992 996 935 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00991 997 996 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00990 1803 1881 996 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00989 935 991 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00988 1803 1000 991 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00987 1087 988 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00986 1803 988 1087 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00985 990 992 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00984 1803 1783 930 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00983 930 1385 929 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00982 929 1034 1059 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00981 1803 1845 938 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00980 938 1087 1003 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00979 1803 931 979 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00978 982 979 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00977 1803 1783 982 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00976 1803 1783 932 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00975 932 1551 986 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00974 984 982 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00973 984 1806 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00972 1803 1385 984 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00971 1803 984 981 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00970 959 962 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00969 922 1845 977 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00968 1803 959 922 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00967 1803 974 926 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00966 926 978 975 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00965 923 971 964 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00964 1803 962 923 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00963 964 972 967 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00962 1803 967 924 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00961 924 972 969 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00960 969 971 925 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00959 972 971 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00958 1803 1881 971 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00957 925 970 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00956 1803 975 970 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00955 962 964 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00954 1803 964 962 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00953 967 969 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00952 1803 977 928 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00951 928 986 927 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00950 927 1150 978 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00949 1803 956 957 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00948 956 962 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00947 1803 921 1033 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00946 919 1031 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00945 920 1218 919 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00944 921 918 920 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00943 912 916 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00942 1803 915 916 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00941 917 1036 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00940 916 914 917 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00939 913 1104 915 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00938 915 918 913 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00937 913 1783 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00936 902 911 904 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00935 1803 918 902 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00934 904 908 903 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00933 1803 903 905 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00932 905 908 909 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00931 909 911 910 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00930 908 911 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00929 1803 1881 911 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00928 910 907 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00927 1803 906 907 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00926 918 904 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00925 1803 904 918 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00924 903 909 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00923 1803 897 899 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00922 899 1217 901 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00921 901 898 900 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00920 900 912 906 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00919 1803 1207 890 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00918 890 889 897 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00917 1803 880 878 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00916 876 1034 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00915 877 1068 876 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00914 880 1035 877 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00913 893 1016 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00912 893 891 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00911 1803 892 893 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00910 1803 893 894 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00909 1803 1783 896 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00908 896 894 895 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00907 895 1101 1020 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00906 887 1035 885 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00905 1803 1034 888 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00904 885 1218 884 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00903 888 1031 887 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00902 1803 884 886 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00901 1803 870 873 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00900 873 874 871 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00899 871 1073 872 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00898 1803 1385 875 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00897 875 889 874 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00896 883 1783 882 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00895 1803 883 889 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00894 882 918 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00893 1803 1385 881 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00892 881 879 999 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00891 1803 867 868 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00890 868 1016 1264 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00889 1803 867 858 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00888 858 891 1241 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00887 1803 1845 857 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00886 857 1399 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00885 857 1385 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00884 859 869 863 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00883 1803 1072 859 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00882 863 866 860 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00881 1803 860 861 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00880 861 866 862 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00879 862 869 865 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00878 866 869 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00877 1803 1881 869 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00876 865 864 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00875 1803 872 864 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00874 1072 863 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00873 1803 863 1072 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00872 860 862 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00871 844 853 843 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00870 1803 841 844 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00869 843 850 842 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00868 1803 842 847 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00867 847 850 848 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00866 848 853 849 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00865 850 853 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00864 1803 1881 853 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00863 849 846 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00862 1803 845 846 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00861 841 843 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00860 1803 843 841 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00859 842 848 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00858 1803 1783 855 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00857 855 854 856 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00856 1803 833 831 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00855 833 841 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00854 1803 834 836 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00853 836 1151 837 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00852 837 1150 839 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00851 835 841 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00850 832 1845 834 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00849 1803 835 832 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00848 1803 977 852 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00847 852 1385 851 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00846 851 856 974 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00845 1803 838 840 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00844 840 839 845 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00843 1803 918 821 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00842 810 812 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00841 1803 813 810 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00840 824 1101 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00839 1803 822 824 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00838 1803 828 824 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00837 824 821 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00836 1803 828 737 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00835 737 826 914 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00834 914 827 736 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00833 736 892 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00832 1803 892 826 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00831 827 828 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00830 1803 1068 723 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00829 723 1035 724 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00828 724 815 725 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00827 725 824 1023 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00826 805 800 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00825 800 1207 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00824 1803 757 800 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00823 1803 892 804 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00822 1803 810 715 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00821 715 759 714 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00820 714 806 898 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00819 822 801 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00818 801 894 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00817 1803 757 801 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00816 815 812 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00815 1803 813 815 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00814 806 918 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00813 1803 805 806 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00812 1803 1029 806 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00811 806 804 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00810 1803 867 752 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00809 752 1029 753 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00808 1803 812 1034 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00807 1803 867 750 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00806 750 804 751 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00805 1803 1218 813 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00804 1803 798 799 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00803 747 981 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00802 748 751 747 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00801 798 796 748 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00800 1803 1845 749 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00799 749 1072 870 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00798 1803 1783 754 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00797 754 813 755 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00796 676 786 788 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00795 1803 931 676 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00794 788 782 789 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00793 1803 789 679 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00792 679 782 787 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00791 787 786 683 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00790 782 786 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00789 1803 1881 786 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00788 683 793 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00787 1803 799 793 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00786 931 788 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00785 1803 788 931 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00784 789 787 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00783 659 764 769 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00782 1803 762 659 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00781 769 763 767 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00780 1803 767 660 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00779 660 763 765 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00778 765 764 663 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00777 763 764 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00776 1803 1881 764 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00775 663 770 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00774 1803 781 770 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00773 762 769 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00772 1803 769 762 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00771 767 765 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00770 796 795 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00769 795 931 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00768 1803 1783 795 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00767 1803 1845 777 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00766 777 1752 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00765 777 1385 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00764 1803 780 781 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00763 744 1252 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00762 745 753 744 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00761 780 774 745 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00760 774 773 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00759 773 762 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00758 1803 1783 773 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00757 1803 834 649 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00756 649 1385 650 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00755 650 755 838 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00754 1803 760 761 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00753 760 931 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00752 711 713 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00751 713 716 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00750 1803 1029 713 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00749 1803 918 718 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00748 718 1029 719 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00747 1803 727 729 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00746 729 728 730 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00745 730 726 738 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00744 731 742 735 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00743 1803 892 731 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00742 735 741 732 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00741 1803 732 733 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00740 733 741 734 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00739 734 742 739 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00738 741 742 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00737 1803 1881 742 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00736 739 740 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00735 1803 738 740 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00734 892 735 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00733 1803 735 892 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00732 732 734 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00731 1803 720 721 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00730 721 804 722 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00729 722 719 728 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00728 700 918 699 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00727 1803 804 696 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00726 699 710 698 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00725 696 1101 700 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00724 1803 698 697 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00723 727 717 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00722 717 716 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00721 1803 804 717 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00720 716 709 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00719 1803 707 709 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00718 708 886 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00717 709 1068 708 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00716 707 706 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00715 706 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00714 1803 1104 706 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00713 1803 710 712 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00712 712 1015 1207 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00711 1803 703 1031 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00710 1803 705 701 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00709 702 1029 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00708 704 1015 702 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00707 705 1218 704 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00706 1803 692 691 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00705 692 703 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00704 1803 867 689 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00703 688 689 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00702 1803 1101 688 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00701 690 695 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00700 1803 691 690 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00699 1803 878 694 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00698 694 701 693 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00697 693 697 695 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00696 687 686 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00695 686 707 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00694 1803 685 686 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00693 668 674 667 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00692 1803 673 668 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00691 667 675 666 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00690 1803 666 670 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00689 670 675 671 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00688 671 674 672 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00687 675 674 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00686 1803 1881 674 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00685 672 669 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00684 1803 678 669 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00683 673 667 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00682 1803 667 673 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00681 666 671 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00680 1803 684 685 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00679 681 867 680 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00678 1803 681 682 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00677 680 685 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00676 1803 682 678 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00675 678 677 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00674 678 857 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00673 1803 648 647 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00672 648 762 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00671 664 661 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00670 1803 1783 664 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00669 654 662 653 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00668 1803 661 654 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00667 653 658 655 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00666 1803 655 651 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00665 651 658 652 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00664 652 662 657 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00663 658 662 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00662 1803 1881 662 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00661 657 656 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00660 1803 665 656 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00659 661 653 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00658 1803 653 661 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00657 655 652 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00656 677 673 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00655 1803 1783 677 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00654 1803 664 665 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00653 665 688 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00652 665 777 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00651 624 622 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00650 559 1029 623 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00649 1803 624 559 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00648 1803 623 549 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00647 549 711 550 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00646 550 616 617 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00645 1803 1207 542 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00644 542 892 543 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00643 543 615 726 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00642 720 619 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00641 1803 1207 720 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00640 622 620 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00639 620 619 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00638 1803 618 620 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00637 1803 891 606 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00636 606 604 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00635 606 892 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00634 1803 710 540 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00633 540 892 538 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00632 538 1015 618 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00631 611 813 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00630 1803 1016 611 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00629 1803 828 611 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00628 611 892 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00627 608 611 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00626 1803 618 547 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00625 547 828 546 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00624 546 615 616 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00623 613 1783 536 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00622 1803 613 879 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00621 536 1035 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00620 519 602 595 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00619 1803 684 519 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00618 595 603 597 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00617 1803 597 522 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00616 522 603 600 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00615 600 602 521 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00614 603 602 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00613 1803 1881 602 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00612 521 601 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00611 1803 596 601 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00610 684 595 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00609 1803 595 684 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00608 597 600 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00607 1803 1101 510 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00606 510 918 592 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00605 593 1783 512 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00604 1803 593 867 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00603 512 1385 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00602 589 583 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00601 1803 588 589 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00600 1803 584 589 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00599 589 684 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00598 1803 590 505 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00597 505 589 507 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00596 507 606 506 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00595 506 1008 591 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00594 579 684 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00593 1803 583 579 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00592 1803 560 576 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00591 497 581 596 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00590 596 687 497 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00589 497 591 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00588 569 1783 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00587 1803 576 569 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00586 1803 569 572 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00585 572 1417 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00584 572 1385 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00583 573 572 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00582 1803 575 573 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00581 493 867 577 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00580 1803 583 493 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00579 494 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00578 577 576 494 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00577 1803 577 575 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00576 1803 564 475 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00575 475 567 563 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00574 1803 565 476 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00573 476 1385 473 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00572 473 566 564 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00571 1803 566 480 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00570 480 1181 481 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00569 481 1150 567 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00568 1803 1385 1150 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00567 562 561 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00566 467 1845 566 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00565 1803 562 467 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00564 1803 1218 539 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00563 539 1015 537 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00562 1803 541 1208 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00561 541 544 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00560 1803 828 1029 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00559 619 545 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00558 545 813 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00557 1803 544 545 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00556 1803 533 535 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00555 535 534 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00554 535 537 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00553 548 558 554 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00552 1803 828 548 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00551 554 557 553 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00550 1803 553 551 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00549 551 557 552 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00548 552 558 555 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00547 557 558 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00546 1803 1881 558 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00545 555 556 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00544 1803 617 556 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00543 828 554 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00542 1803 554 828 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00541 553 552 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00540 1803 531 528 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00539 528 526 529 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00538 529 527 530 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00537 530 535 524 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00536 531 604 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00535 1803 891 531 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00534 1803 828 531 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00533 531 892 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00532 1803 513 518 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00531 518 520 515 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00530 515 514 516 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00529 516 532 517 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00528 1803 891 532 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00527 532 828 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00526 532 892 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00525 1217 509 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00524 509 517 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00523 1803 508 509 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00522 525 1218 523 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00521 1803 525 520 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00520 523 1015 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00519 513 511 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00518 1803 534 513 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00517 1803 918 502 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00516 502 1101 504 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00515 504 854 503 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00514 503 501 508 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00513 1803 579 526 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00512 526 588 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00511 526 495 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00510 499 690 500 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00509 500 498 499 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00508 499 524 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00507 590 534 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00506 1803 592 590 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00505 565 491 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00504 491 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00503 1803 495 491 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00502 1803 495 584 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00501 1803 579 492 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00500 501 492 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00499 1803 565 501 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00498 496 584 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00497 496 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00496 1803 1104 496 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00495 1803 496 498 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00494 1803 466 465 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00493 466 1072 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00492 1803 464 463 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00491 464 673 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00490 483 488 482 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00489 1803 495 483 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00488 482 490 484 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00487 1803 484 487 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00486 487 490 485 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00485 485 488 486 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00484 490 488 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00483 1803 1881 488 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00482 486 489 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00481 1803 500 489 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00480 495 482 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00479 1803 482 495 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00478 484 485 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00477 468 477 469 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00476 1803 560 468 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00475 469 479 470 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00474 1803 470 474 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00473 474 479 471 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00472 471 477 472 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00471 479 477 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00470 1803 1881 477 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00469 472 478 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00468 1803 573 478 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00467 560 469 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00466 1803 469 560 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00465 470 471 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00464 514 812 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00463 1803 419 514 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00462 1803 425 356 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00461 356 424 431 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00460 357 435 427 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00459 1803 1035 357 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00458 427 434 428 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00457 1803 428 362 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00456 362 434 430 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00455 430 435 363 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00454 434 435 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00453 1803 1881 435 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00452 363 432 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00451 1803 431 432 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00450 1035 427 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00449 1803 427 1035 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00448 428 430 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00447 422 420 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00446 422 812 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00445 1803 419 422 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00444 1803 422 424 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00443 1803 1101 351 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00442 351 918 533 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00441 414 396 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00440 343 393 396 1803 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00439 1803 402 343 1803 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00438 343 608 1803 1803 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00437 1803 391 343 1803 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00436 396 400 341 1803 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_00435 341 392 342 1803 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_00434 342 397 1803 1803 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_00433 400 399 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00432 1803 407 400 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00431 393 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00430 1803 583 393 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00429 405 419 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00428 405 812 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00427 1803 511 405 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00426 1803 405 402 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00425 1803 418 420 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00424 1803 695 340 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00423 340 390 392 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00422 348 415 409 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00421 1803 407 348 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00420 409 417 410 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00419 1803 410 350 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00418 350 417 412 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00417 412 415 349 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00416 417 415 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00415 1803 1881 415 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00414 349 416 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00413 1803 414 416 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00412 407 409 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00411 1803 409 407 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00410 410 412 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00409 1803 407 583 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00408 1803 389 339 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00407 339 1101 338 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00406 338 918 337 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00405 337 710 391 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00404 1803 381 322 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00403 322 854 323 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00402 323 390 703 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00401 329 495 328 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00400 1803 390 330 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00399 328 854 384 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00398 330 383 329 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00397 1803 384 389 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00396 386 695 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00395 1803 583 386 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00394 377 380 319 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00393 319 684 377 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00392 1803 390 319 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00391 378 377 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00390 385 389 331 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00389 1803 385 581 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00388 331 386 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00387 1803 382 383 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00386 382 381 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00385 1803 365 364 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 365 661 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00383 1803 1783 317 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 317 374 1382 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 311 375 367 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00380 1803 561 311 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00379 367 373 368 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00378 1803 368 312 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00377 312 373 370 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00376 370 375 316 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00375 373 375 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00374 1803 1881 375 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00373 316 371 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00372 1803 563 371 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00371 561 367 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00370 1803 367 561 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00369 368 370 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00368 1803 1783 318 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00367 318 376 1154 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00366 1803 386 380 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00365 1803 1035 419 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00364 355 1104 354 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00363 354 1035 355 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00362 355 352 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00361 304 359 303 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00360 1803 302 305 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00359 303 354 353 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00358 305 1217 304 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00357 1803 353 425 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00356 358 333 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00355 1803 306 358 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00354 1803 358 361 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00353 361 812 360 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00352 360 419 359 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00351 1803 306 300 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00350 300 879 302 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00349 759 511 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00348 1803 419 759 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00347 347 419 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00346 1803 345 347 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00345 1803 511 347 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00344 347 812 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00343 544 347 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00342 1803 710 891 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00341 1803 419 527 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00340 527 812 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00339 527 511 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00338 344 292 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00337 344 604 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00336 1803 534 344 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00335 1803 344 345 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 1803 346 757 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00333 346 345 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00332 1803 604 854 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00331 1803 334 588 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00330 334 292 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00329 1803 854 418 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00328 418 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00327 418 534 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00326 324 383 326 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00325 1803 324 327 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00324 326 325 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00323 333 332 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00322 332 588 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00321 1803 534 332 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00320 288 534 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00319 287 336 397 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00318 1803 288 287 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00317 335 584 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00316 335 286 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00315 1803 604 335 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00314 1803 335 336 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00313 325 495 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00312 1803 604 325 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00311 1803 1845 1783 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00310 320 327 281 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00309 281 534 320 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00308 1803 279 281 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00307 321 320 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00306 1803 278 275 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00305 275 378 276 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00304 1803 308 309 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 308 561 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00302 268 274 310 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00301 1803 534 268 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00300 310 273 315 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00299 1803 315 314 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00298 314 273 313 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00297 313 274 271 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00296 273 274 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00295 1803 1881 274 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00294 271 272 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00293 1803 321 272 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00292 534 310 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 1803 310 534 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 315 313 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00289 279 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00288 1803 378 279 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00287 615 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00286 1803 534 615 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00285 184 264 260 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00284 1803 812 184 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00283 260 265 257 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00282 1803 257 185 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00281 185 265 259 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00280 259 264 186 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00279 265 264 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00278 1803 1881 264 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00277 186 262 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00276 1803 261 262 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00275 812 260 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 1803 260 812 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00273 257 259 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00272 1803 248 180 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00271 180 250 179 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00270 179 247 261 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00269 254 812 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00268 183 253 255 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 1803 254 183 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00266 1803 306 182 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00265 182 812 181 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00264 181 615 250 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00263 266 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00262 1803 891 266 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00261 1803 244 177 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 177 812 248 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00259 242 399 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00258 1803 710 242 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00257 352 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00256 1803 251 352 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00255 247 245 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00254 1803 255 245 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00253 178 1035 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00252 245 854 178 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00251 175 1035 174 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00250 1803 812 176 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00249 174 1015 240 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00248 176 710 175 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00247 1803 240 241 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00246 172 238 233 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00245 233 757 172 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 172 232 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 234 235 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00242 1803 233 235 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00241 171 418 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00240 235 238 171 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00239 237 511 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00238 173 241 238 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 1803 237 173 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 1803 244 170 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00235 170 604 232 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 1803 383 244 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00233 244 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00232 244 1104 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00231 1803 286 169 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 169 390 231 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 213 376 163 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00228 1803 213 381 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00227 163 211 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00226 1803 190 188 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00225 190 560 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00224 230 383 168 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00223 1803 230 251 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00222 168 390 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00221 227 226 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00220 167 223 292 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 1803 227 167 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 164 224 217 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00217 1803 604 164 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00216 217 225 218 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00215 1803 218 166 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00214 166 225 221 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00213 221 224 165 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00212 225 224 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00211 1803 1881 224 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00210 165 219 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00209 1803 234 219 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00208 604 217 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 1803 217 604 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 218 221 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00205 286 215 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 215 226 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00203 1803 374 215 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00202 1803 202 208 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00201 208 534 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00200 208 212 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00199 1803 1783 162 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 162 276 161 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 161 200 203 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 1803 325 210 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00195 212 210 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00194 1803 226 212 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00193 204 203 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00192 1803 208 204 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00191 158 201 192 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00190 1803 189 158 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00189 192 198 193 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00188 1803 193 159 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00187 159 198 195 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00186 195 201 160 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00185 198 201 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00184 1803 1881 201 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00183 160 197 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00182 1803 204 197 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00181 189 192 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 1803 192 189 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 193 195 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00178 1803 266 156 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00177 156 155 157 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 1803 1217 151 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 151 157 149 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 149 148 150 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 1803 251 154 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00172 154 1015 153 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 153 1068 155 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 253 333 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00169 1803 306 253 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00168 125 124 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 124 122 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00166 1803 534 124 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00165 144 137 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00164 1803 134 137 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00163 136 135 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00162 137 1015 136 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00161 130 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00160 1803 1068 130 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00159 133 131 132 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00158 1803 130 133 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00157 129 352 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00156 132 1068 129 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00155 1803 132 135 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 1803 242 127 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00153 127 231 126 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 126 125 148 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 138 147 139 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00150 1803 1015 138 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00149 139 146 140 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00148 1803 140 141 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00147 141 146 143 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00146 143 147 142 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00145 146 147 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00144 1803 1881 147 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00143 142 145 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00142 1803 144 145 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00141 1015 139 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 1803 139 1015 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 140 143 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00138 111 1068 110 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 1803 111 118 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 110 390 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 121 1015 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00134 121 399 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00133 1803 118 121 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00132 1803 121 117 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00131 109 278 108 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00130 1803 109 112 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 108 226 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 1803 112 113 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00127 113 390 131 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 116 114 134 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 134 117 116 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 116 1217 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00123 1803 96 211 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00122 1803 122 103 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00121 103 333 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 102 376 103 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 103 104 102 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 1803 534 390 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 1803 189 95 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 95 93 96 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 1803 97 278 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 97 211 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00113 84 90 85 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00112 1803 226 84 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00111 85 92 86 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00110 1803 86 87 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00109 87 92 89 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00108 89 90 88 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 92 90 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00106 1803 1881 90 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00105 88 91 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00104 1803 102 91 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00103 226 85 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 1803 85 226 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 86 89 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00100 107 1104 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00099 107 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00098 1803 278 107 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00097 1803 107 104 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 1803 94 202 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 94 96 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00094 1803 226 99 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 99 189 114 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00092 114 534 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 1803 189 374 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 1803 80 18 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 18 79 83 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 83 81 17 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 17 187 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 1803 187 79 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00085 81 80 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00084 1803 122 10 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 10 710 306 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 52 1015 9 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 1803 52 122 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 9 1068 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 14 76 73 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00078 1803 710 14 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00077 73 75 69 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00076 1803 69 16 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00075 16 75 71 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00074 71 76 15 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00073 75 76 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00072 1803 1881 76 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00071 15 74 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00070 1803 150 74 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 710 73 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 1803 73 710 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 69 71 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00066 77 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00065 1803 83 77 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00064 1803 511 1068 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 11 62 55 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00062 1803 53 11 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00061 55 64 57 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00060 1803 57 12 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00059 12 64 59 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00058 59 62 13 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00057 64 62 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 1803 1881 62 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00055 13 63 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 1803 77 63 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00053 53 55 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 1803 55 53 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 57 59 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00050 6 50 43 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00049 1803 511 6 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00048 43 51 44 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 1803 44 8 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 8 51 45 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 45 50 7 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00044 51 50 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00043 1803 1881 50 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00042 7 49 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00041 1803 48 49 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00040 511 43 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 1803 43 511 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 44 45 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00037 48 41 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 1803 38 41 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00035 5 511 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 41 39 5 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 32 80 2 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 1803 32 1104 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 2 534 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 1803 37 38 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 3 34 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 4 226 3 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 37 118 4 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 1803 112 39 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00025 39 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00024 39 1104 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 1803 33 34 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 33 223 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00021 27 53 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 93 27 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 1803 27 93 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 1803 27 93 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 93 27 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 1803 31 399 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 31 30 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00014 1803 28 80 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 28 93 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00012 1803 53 24 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 24 53 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 1803 226 376 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 1803 374 1 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 1 26 200 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 223 374 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 1803 30 223 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 1803 25 26 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 25 24 1803 1803 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00003 30 21 1803 1803 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 21 1845 1803 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 1803 24 21 1803 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C1883 21 1803 1.8635e-14
C1880 24 1803 8.098e-14
C1879 25 1803 1.568e-14
C1878 26 1803 5.238e-14
C1877 27 1803 4.103e-14
C1876 28 1803 1.568e-14
C1874 30 1803 1.3111e-13
C1873 31 1803 1.568e-14
C1872 32 1803 1.8635e-14
C1871 33 1803 1.568e-14
C1870 34 1803 5.023e-14
C1867 37 1803 2.605e-14
C1866 38 1803 7.061e-14
C1865 39 1803 5.343e-14
C1864 40 1803 6.05e-15
C1863 41 1803 1.767e-14
C1861 43 1803 2.871e-14
C1860 44 1803 2.005e-14
C1859 45 1803 2.632e-14
C1856 48 1803 7.038e-14
C1855 49 1803 2.321e-14
C1854 50 1803 5.165e-14
C1853 51 1803 4.869e-14
C1852 52 1803 1.8635e-14
C1851 53 1803 2.5268e-13
C1849 55 1803 2.871e-14
C1848 56 1803 7.43e-15
C1847 57 1803 2.005e-14
C1845 59 1803 2.632e-14
C1843 61 1803 6.05e-15
C1842 62 1803 5.165e-14
C1841 63 1803 2.321e-14
C1840 64 1803 4.869e-14
C1835 69 1803 2.005e-14
C1833 71 1803 2.632e-14
C1831 73 1803 2.871e-14
C1830 74 1803 2.321e-14
C1829 75 1803 4.869e-14
C1828 76 1803 5.165e-14
C1827 77 1803 8.042e-14
C1825 79 1803 2.596e-14
C1824 80 1803 2.4548e-13
C1823 81 1803 2.16e-14
C1822 82 1803 7.76e-15
C1821 83 1803 5.694e-14
C1819 85 1803 2.871e-14
C1818 86 1803 2.005e-14
C1815 89 1803 2.632e-14
C1814 90 1803 5.165e-14
C1813 91 1803 2.321e-14
C1812 92 1803 4.869e-14
C1811 93 1803 1.1467e-13
C1810 94 1803 1.568e-14
C1808 96 1803 8.306e-14
C1807 97 1803 1.568e-14
C1806 98 1803 6.05e-15
C1802 102 1803 9.738e-14
C1801 103 1803 7.43e-15
C1800 104 1803 4.487e-14
C1797 107 1803 2.455e-14
C1795 109 1803 1.8635e-14
C1793 111 1803 1.8635e-14
C1792 112 1803 1.0177e-13
C1790 114 1803 1.0909e-13
C1788 116 1803 4.11e-15
C1787 117 1803 4.997e-14
C1786 118 1803 1.0352e-13
C1783 121 1803 2.455e-14
C1782 122 1803 2.098e-13
C1780 124 1803 1.8635e-14
C1779 125 1803 5.396e-14
C1774 130 1803 5.521e-14
C1773 131 1803 9.921e-14
C1772 132 1803 2.445e-14
C1770 134 1803 1.0213e-13
C1769 135 1803 5.833e-14
C1767 137 1803 1.767e-14
C1765 139 1803 2.871e-14
C1764 140 1803 2.005e-14
C1761 143 1803 2.632e-14
C1760 144 1803 6.918e-14
C1759 145 1803 2.321e-14
C1758 146 1803 4.869e-14
C1757 147 1803 5.165e-14
C1756 148 1803 1.116e-13
C1754 150 1803 5.626e-14
C1749 155 1803 5.75e-14
C1746 157 1803 7.006e-14
C1731 172 1803 4.11e-15
C1716 187 1803 6.68e-14
C1714 188 1803 2.899e-14
C1713 189 1803 1.6583e-13
C1712 190 1803 1.568e-14
C1710 192 1803 2.871e-14
C1709 193 1803 2.005e-14
C1707 195 1803 2.632e-14
C1705 197 1803 2.321e-14
C1704 198 1803 4.869e-14
C1702 200 1803 6.546e-14
C1701 201 1803 5.165e-14
C1700 202 1803 5.608e-14
C1699 203 1803 5.49e-14
C1698 204 1803 6.002e-14
C1694 208 1803 5.422e-14
C1692 210 1803 1.677e-14
C1691 211 1803 9.566e-14
C1690 212 1803 5.188e-14
C1689 213 1803 1.8635e-14
C1687 215 1803 1.8635e-14
C1685 217 1803 2.871e-14
C1684 218 1803 2.005e-14
C1683 219 1803 2.321e-14
C1681 221 1803 2.632e-14
C1679 223 1803 1.1619e-13
C1678 224 1803 5.165e-14
C1677 225 1803 4.869e-14
C1676 226 1803 3.59e-13
C1675 227 1803 1.662e-14
C1672 230 1803 1.8635e-14
C1671 231 1803 9.286e-14
C1670 232 1803 5.121e-14
C1669 233 1803 5.293e-14
C1668 234 1803 8.838e-14
C1667 235 1803 1.767e-14
C1665 237 1803 1.662e-14
C1664 238 1803 6.948e-14
C1663 239 1803 6.05e-15
C1662 240 1803 2.306e-14
C1661 241 1803 5.51e-14
C1660 242 1803 5.871e-14
C1658 244 1803 1.4138e-13
C1657 245 1803 1.767e-14
C1656 246 1803 6.05e-15
C1655 247 1803 5.852e-14
C1654 248 1803 6.521e-14
C1652 250 1803 6.34e-14
C1651 251 1803 2.1493e-13
C1649 253 1803 7.566e-14
C1648 254 1803 1.662e-14
C1647 255 1803 8.687e-14
C1645 257 1803 2.005e-14
C1643 259 1803 2.632e-14
C1642 260 1803 2.871e-14
C1641 261 1803 9.826e-14
C1640 262 1803 2.321e-14
C1638 264 1803 5.165e-14
C1637 265 1803 4.869e-14
C1636 266 1803 5.433e-14
C1630 272 1803 2.321e-14
C1629 273 1803 4.869e-14
C1628 274 1803 5.165e-14
C1626 276 1803 6.286e-14
C1624 278 1803 1.6321e-13
C1623 279 1803 5.397e-14
C1621 281 1803 4.11e-15
C1616 286 1803 1.265e-13
C1614 288 1803 1.662e-14
C1610 292 1803 1.3514e-13
C1600 302 1803 6.756e-14
C1596 306 1803 2.3326e-13
C1593 308 1803 1.568e-14
C1592 309 1803 3.067e-14
C1591 310 1803 2.871e-14
C1588 313 1803 2.632e-14
C1586 315 1803 2.005e-14
C1582 319 1803 4.11e-15
C1581 320 1803 1.853e-14
C1580 321 1803 7.038e-14
C1577 324 1803 1.8635e-14
C1576 325 1803 1.0882e-13
C1574 327 1803 4.513e-14
C1569 332 1803 1.8635e-14
C1568 333 1803 2.8696e-13
C1567 334 1803 1.568e-14
C1566 335 1803 2.455e-14
C1565 336 1803 7.042e-14
C1558 343 1803 4.11e-15
C1557 344 1803 2.455e-14
C1556 345 1803 9.932e-14
C1555 346 1803 1.568e-14
C1554 347 1803 2.72e-14
C1549 352 1803 1.2032e-13
C1548 353 1803 2.306e-14
C1547 354 1803 5.147e-14
C1546 355 1803 4.11e-15
C1543 358 1803 5.751e-14
C1542 359 1803 6.15e-14
C1536 364 1803 2.371e-14
C1535 365 1803 1.568e-14
C1533 367 1803 2.871e-14
C1532 368 1803 2.005e-14
C1530 370 1803 2.632e-14
C1529 371 1803 2.321e-14
C1527 373 1803 4.869e-14
C1526 374 1803 2.2494e-13
C1525 375 1803 5.165e-14
C1524 376 1803 2.0442e-13
C1523 377 1803 1.853e-14
C1522 378 1803 8.936e-14
C1520 380 1803 4.329e-14
C1519 381 1803 1.0716e-13
C1518 382 1803 1.568e-14
C1517 383 1803 1.7618e-13
C1516 384 1803 2.306e-14
C1515 385 1803 1.8635e-14
C1514 386 1803 1.2612e-13
C1511 389 1803 1.0227e-13
C1510 390 1803 3.7963e-13
C1509 391 1803 6.647e-14
C1508 392 1803 5.361e-14
C1507 393 1803 7.306e-14
C1504 396 1803 2.259e-14
C1503 397 1803 5.469e-14
C1502 398 1803 9.96e-15
C1501 399 1803 2.2065e-13
C1500 400 1803 5.056e-14
C1498 402 1803 7.127e-14
C1495 405 1803 2.455e-14
C1493 407 1803 1.5659e-13
C1491 409 1803 2.871e-14
C1490 410 1803 2.005e-14
C1488 412 1803 2.632e-14
C1486 414 1803 8.594e-14
C1485 415 1803 5.165e-14
C1484 416 1803 2.321e-14
C1483 417 1803 4.869e-14
C1482 418 1803 1.5916e-13
C1481 419 1803 2.9519e-13
C1480 420 1803 5.019e-14
C1478 422 1803 2.455e-14
C1476 424 1803 5.842e-14
C1475 425 1803 6.305e-14
C1473 427 1803 2.871e-14
C1472 428 1803 2.005e-14
C1470 430 1803 2.632e-14
C1469 431 1803 6.412e-14
C1468 432 1803 2.321e-14
C1466 434 1803 4.869e-14
C1465 435 1803 5.165e-14
C1436 463 1803 8.683e-14
C1435 464 1803 1.568e-14
C1434 465 1803 2.899e-14
C1433 466 1803 1.568e-14
C1430 469 1803 2.871e-14
C1429 470 1803 2.005e-14
C1428 471 1803 2.632e-14
C1422 477 1803 5.165e-14
C1421 478 1803 2.321e-14
C1420 479 1803 4.869e-14
C1417 482 1803 2.871e-14
C1415 484 1803 2.005e-14
C1414 485 1803 2.632e-14
C1411 488 1803 5.165e-14
C1410 489 1803 2.321e-14
C1409 490 1803 4.869e-14
C1408 491 1803 1.8635e-14
C1407 492 1803 1.677e-14
C1404 495 1803 2.1548e-13
C1403 496 1803 2.455e-14
C1402 497 1803 4.11e-15
C1401 498 1803 5.597e-14
C1400 499 1803 4.11e-15
C1399 500 1803 8.418e-14
C1398 501 1803 8.89e-14
C1391 508 1803 6.221e-14
C1390 509 1803 1.8635e-14
C1388 511 1803 4.0353e-13
C1386 513 1803 5.416e-14
C1385 514 1803 6.676e-14
C1382 517 1803 6.497e-14
C1379 520 1803 4.978e-14
C1375 524 1803 1.0631e-13
C1374 525 1803 1.8635e-14
C1373 526 1803 1.3498e-13
C1372 527 1803 7.132e-14
C1368 531 1803 5.836e-14
C1367 532 1803 8.992e-14
C1366 533 1803 5.826e-14
C1365 534 1803 7.53399e-13
C1364 535 1803 8.032e-14
C1362 537 1803 5.076e-14
C1358 541 1803 1.568e-14
C1355 544 1803 1.3738e-13
C1354 545 1803 1.8635e-14
C1347 552 1803 2.632e-14
C1346 553 1803 2.005e-14
C1345 554 1803 2.871e-14
C1343 556 1803 2.321e-14
C1342 557 1803 4.869e-14
C1341 558 1803 5.165e-14
C1338 560 1803 1.4314e-13
C1337 561 1803 1.27e-13
C1336 562 1803 1.662e-14
C1335 563 1803 6.412e-14
C1334 564 1803 5.225e-14
C1333 565 1803 1.1747e-13
C1332 566 1803 9.417e-14
C1331 567 1803 5.99e-14
C1329 569 1803 5.056e-14
C1326 572 1803 5.482e-14
C1325 573 1803 8.162e-14
C1323 575 1803 4.798e-14
C1322 576 1803 1.3005e-13
C1321 577 1803 2.445e-14
C1320 578 1803 7.43e-15
C1319 579 1803 9.409e-14
C1317 581 1803 7.531e-14
C1315 583 1803 2.0327e-13
C1314 584 1803 1.43e-13
C1310 588 1803 1.5768e-13
C1309 589 1803 5.806e-14
C1308 590 1803 5.416e-14
C1307 591 1803 6.791e-14
C1306 592 1803 5.616e-14
C1305 593 1803 1.8635e-14
C1303 595 1803 2.871e-14
C1302 596 1803 9.858e-14
C1301 597 1803 2.005e-14
C1298 600 1803 2.632e-14
C1297 601 1803 2.321e-14
C1296 602 1803 5.165e-14
C1295 603 1803 4.869e-14
C1294 604 1803 3.5668e-13
C1292 606 1803 1.0012e-13
C1290 608 1803 1.0357e-13
C1287 611 1803 2.72e-14
C1285 613 1803 1.8635e-14
C1283 615 1803 1.6296e-13
C1282 616 1803 5.76e-14
C1281 617 1803 6.826e-14
C1280 618 1803 1.1436e-13
C1279 619 1803 1.0743e-13
C1278 620 1803 1.8635e-14
C1276 622 1803 5.785e-14
C1275 623 1803 6.281e-14
C1274 624 1803 1.662e-14
C1257 641 1803 6.05e-15
C1250 647 1803 3.139e-14
C1249 648 1803 1.568e-14
C1245 652 1803 2.632e-14
C1244 653 1803 2.871e-14
C1242 655 1803 2.005e-14
C1241 656 1803 2.321e-14
C1239 658 1803 4.869e-14
C1236 661 1803 1.4321e-13
C1235 662 1803 5.165e-14
C1233 664 1803 4.816e-14
C1232 665 1803 6.338e-14
C1231 666 1803 2.005e-14
C1230 667 1803 2.871e-14
C1228 669 1803 2.321e-14
C1226 671 1803 2.632e-14
C1224 673 1803 1.6433e-13
C1223 674 1803 5.165e-14
C1222 675 1803 4.869e-14
C1220 677 1803 4.981e-14
C1219 678 1803 6.338e-14
C1216 681 1803 1.8635e-14
C1215 682 1803 4.768e-14
C1213 684 1803 2.6504e-13
C1212 685 1803 8.646e-14
C1211 686 1803 1.8635e-14
C1210 687 1803 5.021e-14
C1209 688 1803 1.0783e-13
C1208 689 1803 1.677e-14
C1207 690 1803 6.979e-14
C1206 691 1803 4.798e-14
C1205 692 1803 1.568e-14
C1202 695 1803 1.9221e-13
C1200 697 1803 5.52e-14
C1199 698 1803 2.306e-14
C1196 701 1803 6.7e-14
C1194 703 1803 1.9856e-13
C1192 705 1803 2.605e-14
C1191 706 1803 1.8635e-14
C1190 707 1803 1.4354e-13
C1188 709 1803 1.767e-14
C1187 710 1803 5.0232e-13
C1186 711 1803 9.936e-14
C1184 713 1803 1.8635e-14
C1181 716 1803 1.011e-13
C1180 717 1803 1.8635e-14
C1178 719 1803 5.226e-14
C1177 720 1803 5.751e-14
C1171 726 1803 7.44e-14
C1170 727 1803 7.531e-14
C1169 728 1803 6.1e-14
C1165 732 1803 2.005e-14
C1163 734 1803 2.632e-14
C1162 735 1803 2.871e-14
C1159 738 1803 6.826e-14
C1157 740 1803 2.321e-14
C1156 741 1803 4.869e-14
C1155 742 1803 5.165e-14
C1146 751 1803 5.511e-14
C1144 753 1803 1.0311e-13
C1142 755 1803 1.701e-13
C1140 757 1803 1.9899e-13
C1138 759 1803 1.0436e-13
C1136 760 1803 1.568e-14
C1135 761 1803 2.899e-14
C1134 762 1803 1.2992e-13
C1133 763 1803 4.869e-14
C1132 764 1803 5.165e-14
C1131 765 1803 2.632e-14
C1129 767 1803 2.005e-14
C1127 769 1803 2.871e-14
C1126 770 1803 2.321e-14
C1123 773 1803 1.8635e-14
C1122 774 1803 5.591e-14
C1119 777 1803 6.682e-14
C1116 780 1803 2.605e-14
C1115 781 1803 6.586e-14
C1114 782 1803 4.869e-14
C1110 786 1803 5.165e-14
C1109 787 1803 2.632e-14
C1108 788 1803 2.871e-14
C1107 789 1803 2.005e-14
C1103 793 1803 2.321e-14
C1101 795 1803 1.8635e-14
C1100 796 1803 5.231e-14
C1098 798 1803 2.605e-14
C1097 799 1803 6.346e-14
C1096 800 1803 1.8635e-14
C1095 801 1803 1.8635e-14
C1092 804 1803 2.5969e-13
C1091 805 1803 6.326e-14
C1090 806 1803 5.596e-14
C1086 810 1803 5.631e-14
C1084 812 1803 6.3644e-13
C1083 813 1803 2.907e-13
C1081 815 1803 5.356e-14
C1075 821 1803 6.384e-14
C1074 822 1803 9.686e-14
C1072 824 1803 6.436e-14
C1070 826 1803 2.596e-14
C1069 827 1803 2.16e-14
C1068 828 1803 3.4382e-13
C1067 829 1803 7.76e-15
C1066 830 1803 6.05e-15
C1064 831 1803 2.659e-14
C1062 833 1803 1.568e-14
C1061 834 1803 9.032e-14
C1060 835 1803 1.662e-14
C1057 838 1803 7.265e-14
C1056 839 1803 5.51e-14
C1054 841 1803 1.0972e-13
C1053 842 1803 2.005e-14
C1052 843 1803 2.871e-14
C1050 845 1803 6.172e-14
C1049 846 1803 2.321e-14
C1047 848 1803 2.632e-14
C1045 850 1803 4.869e-14
C1042 853 1803 5.165e-14
C1041 854 1803 3.8296e-13
C1039 856 1803 5.106e-14
C1038 857 1803 7.882e-14
C1035 860 1803 2.005e-14
C1033 862 1803 2.632e-14
C1032 863 1803 2.871e-14
C1031 864 1803 2.321e-14
C1029 866 1803 4.869e-14
C1028 867 1803 3.3727e-13
C1026 869 1803 5.165e-14
C1025 870 1803 5.681e-14
C1023 872 1803 6.106e-14
C1021 874 1803 5.446e-14
C1017 878 1803 7.415e-14
C1016 879 1803 2.0388e-13
C1015 880 1803 2.605e-14
C1012 883 1803 1.8635e-14
C1011 884 1803 2.306e-14
C1009 886 1803 8.625e-14
C1006 889 1803 1.1124e-13
C1004 891 1803 4.8499e-13
C1003 892 1803 4.272e-13
C1002 893 1803 2.455e-14
C1001 894 1803 1.0249e-13
C998 897 1803 7.266e-14
C997 898 1803 5.82e-14
C992 903 1803 2.005e-14
C991 904 1803 2.871e-14
C989 906 1803 7.122e-14
C988 907 1803 2.321e-14
C987 908 1803 4.869e-14
C986 909 1803 2.632e-14
C984 911 1803 5.165e-14
C983 912 1803 9.092e-14
C982 913 1803 4.11e-15
C981 914 1803 5.375e-14
C980 915 1803 5.533e-14
C979 916 1803 1.767e-14
C977 918 1803 5.8237e-13
C974 921 1803 2.605e-14
C964 931 1803 2.1905e-13
C938 956 1803 1.568e-14
C937 957 1803 2.827e-14
C935 959 1803 1.662e-14
C932 962 1803 1.0372e-13
C930 964 1803 2.871e-14
C927 967 1803 2.005e-14
C925 969 1803 2.632e-14
C924 970 1803 2.321e-14
C923 971 1803 5.165e-14
C922 972 1803 4.869e-14
C920 974 1803 5.825e-14
C919 975 1803 5.452e-14
C917 977 1803 1.2944e-13
C916 978 1803 5.63e-14
C915 979 1803 1.677e-14
C913 981 1803 8.195e-14
C912 982 1803 5.053e-14
C910 984 1803 2.455e-14
C908 986 1803 8.086e-14
C906 988 1803 2.871e-14
C904 990 1803 2.005e-14
C903 991 1803 2.321e-14
C902 992 1803 2.632e-14
C898 996 1803 5.165e-14
C897 997 1803 4.869e-14
C895 999 1803 5.566e-14
C894 1000 1803 5.626e-14
C891 1003 1803 5.441e-14
C890 1004 1803 1.8635e-14
C888 1006 1803 5.143e-14
C887 1007 1803 2.605e-14
C886 1008 1803 1.38e-13
C883 1011 1803 1.8635e-14
C882 1012 1803 4.363e-14
C881 1013 1803 5.413e-14
C879 1015 1803 6.7294e-13
C878 1016 1803 2.1844e-13
C877 1017 1803 1.8635e-14
C874 1020 1803 6.491e-14
C873 1021 1803 1.8635e-14
C871 1023 1803 7.976e-14
C868 1026 1803 5.943e-14
C867 1027 1803 5.62e-14
C865 1029 1803 4.5539e-13
C864 1030 1803 5.586e-14
C863 1031 1803 2.2037e-13
C861 1033 1803 5.73e-14
C860 1034 1803 3.811e-13
C859 1035 1803 6.6186e-13
C858 1036 1803 9.546e-14
C857 1037 1803 2.306e-14
C855 1038 1803 7.76e-15
C853 1040 1803 2.871e-14
C852 1041 1803 2.005e-14
C851 1042 1803 2.321e-14
C850 1043 1803 2.632e-14
C847 1046 1803 4.869e-14
C846 1047 1803 5.165e-14
C845 1048 1803 1.8635e-14
C844 1049 1803 5.986e-14
C842 1051 1803 4.991e-14
C841 1052 1803 4.907e-14
C839 1054 1803 2.605e-14
C838 1055 1803 2.455e-14
C837 1056 1803 7.027e-14
C836 1057 1803 1.568e-14
C834 1059 1803 8.085e-14
C833 1060 1803 1.662e-14
C829 1064 1803 6.065e-14
C828 1065 1803 5.63e-14
C826 1067 1803 1.0744e-13
C825 1068 1803 8.19869e-13
C824 1069 1803 5.346e-14
C821 1072 1803 2.8775e-13
C820 1073 1803 7.532e-14
C819 1074 1803 5.011e-14
C818 1075 1803 9.816e-14
C817 1076 1803 2.455e-14
C816 1077 1803 1.8635e-14
C814 1079 1803 2.005e-14
C813 1080 1803 2.871e-14
C812 1081 1803 2.321e-14
C809 1084 1803 2.632e-14
C808 1085 1803 4.869e-14
C807 1086 1803 5.165e-14
C806 1087 1803 2.4583e-13
C805 1088 1803 9.98e-14
C804 1089 1803 5.011e-14
C803 1090 1803 2.455e-14
C801 1092 1803 2.871e-14
C800 1093 1803 2.005e-14
C798 1095 1803 2.632e-14
C796 1097 1803 5.746e-14
C795 1098 1803 5.165e-14
C794 1099 1803 2.321e-14
C793 1100 1803 4.869e-14
C792 1101 1803 5.7109e-13
C791 1102 1803 1.8635e-14
C790 1103 1803 5.856e-14
C789 1104 1803 6.0121e-13
C788 1105 1803 5.926e-14
C787 1106 1803 1.853e-14
C785 1108 1803 4.11e-15
C784 1109 1803 6.157e-14
C783 1110 1803 2.596e-14
C782 1111 1803 9.392e-14
C781 1112 1803 2.16e-14
C762 1131 1803 4.11e-15
C745 1147 1803 1.568e-14
C744 1148 1803 2.371e-14
C743 1149 1803 1.1624e-13
C742 1150 1803 3.1024e-13
C741 1151 1803 8.206e-14
C740 1152 1803 1.662e-14
C738 1154 1803 1.4586e-13
C737 1155 1803 9.277e-14
C736 1156 1803 6.11e-14
C735 1157 1803 5.825e-14
C733 1159 1803 2.871e-14
C732 1160 1803 2.005e-14
C730 1162 1803 2.632e-14
C728 1164 1803 6.172e-14
C727 1165 1803 5.165e-14
C726 1166 1803 2.321e-14
C725 1167 1803 4.869e-14
C724 1168 1803 1.568e-14
C723 1169 1803 1.102e-13
C722 1170 1803 2.005e-14
C720 1172 1803 2.871e-14
C717 1175 1803 5.692e-14
C716 1176 1803 2.321e-14
C714 1178 1803 2.632e-14
C713 1179 1803 4.869e-14
C711 1181 1803 1.6944e-13
C710 1182 1803 5.165e-14
C709 1183 1803 1.8635e-14
C708 1184 1803 5.326e-14
C707 1185 1803 5.655e-14
C705 1187 1803 9.126e-14
C704 1188 1803 4.937e-14
C701 1191 1803 1.767e-14
C700 1192 1803 6.05e-15
C699 1193 1803 6.789e-14
C698 1194 1803 1.1503e-13
C697 1195 1803 8.5e-14
C696 1196 1803 2.306e-14
C695 1197 1803 2.005e-14
C694 1198 1803 2.871e-14
C692 1200 1803 2.321e-14
C690 1202 1803 2.632e-14
C689 1203 1803 4.869e-14
C687 1205 1803 5.165e-14
C686 1206 1803 2.605e-14
C685 1207 1803 3.2507e-13
C684 1208 1803 1.2586e-13
C680 1212 1803 6.51e-14
C679 1213 1803 5.482e-14
C677 1215 1803 5.516e-14
C676 1216 1803 6.546e-14
C675 1217 1803 5.1152e-13
C674 1218 1803 5.3799e-13
C671 1221 1803 2.005e-14
C669 1223 1803 2.632e-14
C668 1224 1803 2.871e-14
C667 1225 1803 6.826e-14
C665 1227 1803 5.165e-14
C664 1228 1803 2.321e-14
C663 1229 1803 4.869e-14
C662 1230 1803 2.371e-14
C657 1235 1803 2.321e-14
C656 1236 1803 4.869e-14
C653 1239 1803 5.165e-14
C652 1240 1803 4.991e-14
C651 1241 1803 1.1031e-13
C648 1244 1803 5.986e-14
C647 1245 1803 1.5449e-13
C645 1247 1803 5.507e-14
C644 1248 1803 1.677e-14
C643 1249 1803 4.813e-14
C640 1252 1803 1.0547e-13
C634 1258 1803 2.321e-14
C630 1262 1803 4.869e-14
C629 1263 1803 5.165e-14
C628 1264 1803 8.871e-14
C625 1267 1803 5.986e-14
C624 1268 1803 4.991e-14
C621 1271 1803 4.907e-14
C618 1274 1803 8.518e-14
C611 1281 1803 7.041e-14
C609 1283 1803 5.39e-14
C605 1287 1803 6.554e-14
C604 1288 1803 6.291e-14
C603 1289 1803 7.43e-15
C597 1295 1803 5.611e-14
C594 1298 1803 4.179e-14
C589 1303 1803 2.321e-14
C588 1304 1803 4.869e-14
C586 1306 1803 8.454e-14
C584 1308 1803 5.165e-14
C579 1313 1803 6.362e-14
C577 1314 1803 2.321e-14
C576 1315 1803 4.869e-14
C575 1316 1803 5.165e-14
C573 1318 1803 1.568e-14
C572 1319 1803 2.871e-14
C570 1321 1803 2.005e-14
C569 1322 1803 2.632e-14
C565 1326 1803 1.8635e-14
C562 1329 1803 2.605e-14
C561 1330 1803 2.455e-14
C560 1331 1803 4.11e-15
C558 1333 1803 2.455e-14
C557 1334 1803 2.871e-14
C556 1335 1803 2.005e-14
C555 1336 1803 2.632e-14
C553 1338 1803 1.8635e-14
C552 1339 1803 4.11e-15
C550 1341 1803 2.605e-14
C548 1343 1803 2.455e-14
C544 1347 1803 2.72e-14
C541 1350 1803 2.72e-14
C538 1353 1803 5.223e-14
C537 1354 1803 6.092e-14
C536 1355 1803 5.88e-14
C533 1358 1803 1.8635e-14
C532 1359 1803 2.445e-14
C531 1360 1803 2.455e-14
C530 1361 1803 2.871e-14
C529 1362 1803 7.43e-15
C528 1363 1803 2.005e-14
C527 1364 1803 2.632e-14
C524 1367 1803 2.871e-14
C522 1369 1803 2.005e-14
C521 1370 1803 2.632e-14
C516 1374 1803 2.871e-14
C515 1375 1803 2.005e-14
C514 1376 1803 2.321e-14
C512 1378 1803 2.632e-14
C510 1380 1803 4.869e-14
C509 1381 1803 5.165e-14
C508 1382 1803 1.6146e-13
C507 1383 1803 1.662e-14
C506 1384 1803 5.655e-14
C505 1385 1803 1.17243e-12
C503 1387 1803 6.378e-14
C502 1388 1803 9.047e-14
C501 1389 1803 1.662e-14
C500 1390 1803 4.611e-14
C499 1391 1803 1.2944e-13
C498 1392 1803 1.568e-14
C496 1394 1803 7.675e-14
C495 1395 1803 5.613e-14
C493 1397 1803 6.05e-15
C492 1398 1803 1.767e-14
C491 1399 1803 3.016e-13
C487 1403 1803 2.72e-14
C485 1405 1803 5.297e-14
C484 1406 1803 5.535e-14
C483 1407 1803 6.963e-14
C482 1408 1803 9.945e-14
C481 1409 1803 2.605e-14
C480 1410 1803 5.475e-14
C479 1411 1803 2.0575e-13
C475 1415 1803 2.605e-14
C474 1416 1803 5.611e-14
C473 1417 1803 3.7214e-13
C471 1419 1803 2.005e-14
C470 1420 1803 2.871e-14
C469 1421 1803 1.2198e-13
C468 1422 1803 4.869e-14
C467 1423 1803 2.321e-14
C465 1425 1803 2.632e-14
C463 1427 1803 5.165e-14
C458 1432 1803 5.449e-14
C457 1433 1803 2.8063e-13
C456 1434 1803 1.8635e-14
C454 1436 1803 7.407e-14
C449 1441 1803 1.506e-13
C447 1443 1803 6.493e-14
C446 1444 1803 5.581e-14
C445 1445 1803 1.767e-14
C444 1446 1803 6.05e-15
C443 1447 1803 1.8635e-14
C442 1448 1803 2.4383e-13
C440 1450 1803 2.871e-14
C439 1451 1803 2.005e-14
C437 1453 1803 2.632e-14
C436 1454 1803 7.758e-14
C435 1455 1803 2.321e-14
C433 1457 1803 5.165e-14
C432 1458 1803 4.869e-14
C424 1466 1803 4.11e-15
C422 1468 1803 8.58e-15
C421 1469 1803 4.209e-14
C420 1470 1803 5.086e-14
C410 1480 1803 5.806e-14
C408 1482 1803 5.461e-14
C401 1489 1803 6.05e-15
C382 1507 1803 1.2115e-13
C381 1508 1803 2.871e-14
C380 1509 1803 2.632e-14
C379 1510 1803 2.005e-14
C378 1511 1803 4.869e-14
C377 1512 1803 2.321e-14
C376 1513 1803 5.05e-14
C372 1517 1803 5.165e-14
C371 1518 1803 2.299e-14
C368 1521 1803 1.8635e-14
C367 1522 1803 7.577e-14
C366 1523 1803 1.8635e-14
C365 1524 1803 8.233e-14
C362 1527 1803 5.367e-14
C357 1532 1803 2.455e-14
C356 1533 1803 4.531e-14
C355 1534 1803 7.585e-14
C354 1535 1803 5.196e-14
C350 1539 1803 1.8635e-14
C349 1540 1803 1.7305e-13
C347 1542 1803 1.8635e-14
C342 1547 1803 2.306e-14
C341 1548 1803 1.0106e-13
C340 1549 1803 1.8635e-14
C338 1551 1803 2.7426e-13
C336 1553 1803 1.3113e-13
C335 1554 1803 7.43e-15
C332 1557 1803 5.041e-14
C330 1559 1803 4.747e-14
C328 1561 1803 3.3546e-13
C327 1562 1803 2.306e-14
C326 1563 1803 1.2873e-13
C323 1566 1803 2.605e-14
C322 1567 1803 1.0174e-13
C319 1570 1803 2.871e-14
C318 1571 1803 2.632e-14
C317 1572 1803 4.11e-15
C316 1573 1803 2.321e-14
C315 1574 1803 1.101e-13
C314 1575 1803 2.005e-14
C313 1576 1803 4.869e-14
C310 1579 1803 5.165e-14
C308 1581 1803 4.11e-15
C305 1584 1803 2.871e-14
C303 1586 1803 2.632e-14
C302 1587 1803 4.869e-14
C300 1589 1803 2.005e-14
C298 1591 1803 2.321e-14
C297 1592 1803 6.378e-14
C296 1593 1803 5.165e-14
C293 1595 1803 1.3012e-13
C292 1596 1803 1.7068e-13
C291 1597 1803 1.568e-14
C290 1598 1803 1.568e-14
C289 1599 1803 2.596e-14
C288 1600 1803 7.76e-15
C287 1601 1803 4.974e-14
C286 1602 1803 2.16e-14
C284 1604 1803 4.786e-14
C283 1605 1803 2.596e-14
C282 1606 1803 2.16e-14
C281 1607 1803 9.7e-15
C280 1608 1803 2.605e-14
C279 1609 1803 2.306e-14
C278 1610 1803 7.854e-14
C277 1611 1803 1.0126e-13
C276 1612 1803 2.605e-14
C275 1613 1803 2.5805e-13
C274 1614 1803 1.662e-14
C273 1615 1803 5.331e-14
C272 1616 1803 6.551e-14
C271 1617 1803 1.767e-14
C270 1618 1803 6.05e-15
C269 1619 1803 1.4885e-13
C268 1620 1803 4.2043e-13
C266 1622 1803 2.605e-14
C265 1623 1803 8.421e-14
C264 1624 1803 1.3712e-13
C263 1625 1803 6.05e-15
C262 1626 1803 2.0416e-13
C261 1627 1803 8.346e-14
C260 1628 1803 2.306e-14
C259 1629 1803 5.727e-14
C258 1630 1803 9.951e-14
C257 1631 1803 2.605e-14
C255 1633 1803 1.8635e-14
C254 1634 1803 6.735e-14
C253 1635 1803 5.231e-14
C251 1637 1803 2.596e-14
C250 1638 1803 9.7e-15
C249 1639 1803 5.215e-14
C248 1640 1803 2.16e-14
C247 1641 1803 5.607e-14
C246 1642 1803 4.4574e-13
C244 1644 1803 2.871e-14
C243 1645 1803 2.005e-14
C242 1646 1803 2.632e-14
C240 1648 1803 8.538e-14
C239 1649 1803 2.321e-14
C237 1651 1803 4.869e-14
C236 1652 1803 5.165e-14
C235 1653 1803 3.547e-14
C230 1658 1803 6.05e-15
C227 1661 1803 8.58e-15
C217 1671 1803 8.58e-15
C213 1675 1803 8.58e-15
C206 1682 1803 6.05e-15
C205 1683 1803 9.7e-15
C202 1685 1803 2.871e-14
C200 1687 1803 2.005e-14
C199 1688 1803 2.321e-14
C197 1690 1803 2.632e-14
C194 1693 1803 4.869e-14
C193 1694 1803 5.165e-14
C191 1696 1803 5.981e-14
C188 1699 1803 2.605e-14
C187 1700 1803 6.078e-14
C185 1702 1803 1.464e-13
C184 1703 1803 5.3621e-13
C182 1705 1803 1.767e-14
C181 1706 1803 4.11e-15
C180 1707 1803 2.605e-14
C175 1712 1803 5.13e-14
C174 1713 1803 6.03e-14
C173 1714 1803 5.041e-14
C172 1715 1803 8.086e-14
C171 1716 1803 2.299e-14
C170 1717 1803 4.11e-15
C168 1719 1803 3.0676e-13
C165 1722 1803 2.005e-14
C163 1724 1803 2.632e-14
C162 1725 1803 2.871e-14
C159 1728 1803 6.85e-14
C158 1729 1803 2.321e-14
C157 1730 1803 4.869e-14
C155 1732 1803 1.7076e-13
C154 1733 1803 1.0193e-13
C153 1734 1803 5.165e-14
C152 1735 1803 7.43e-15
C151 1736 1803 2.5033e-13
C150 1737 1803 8.536e-14
C149 1738 1803 1.677e-14
C147 1740 1803 2.005e-14
C145 1742 1803 2.871e-14
C144 1743 1803 4.869e-14
C143 1744 1803 2.321e-14
C142 1745 1803 2.632e-14
C139 1748 1803 5.165e-14
C138 1749 1803 5.05e-14
C137 1750 1803 6.628e-14
C136 1751 1803 5.454e-14
C135 1752 1803 5.1271e-13
C134 1753 1803 2.299e-14
C133 1754 1803 4.11e-15
C131 1756 1803 4.561e-14
C130 1757 1803 8.02e-14
C129 1758 1803 9.798e-14
C127 1760 1803 2.299e-14
C126 1761 1803 4.11e-15
C124 1763 1803 2.4198e-13
C122 1765 1803 2.005e-14
C120 1767 1803 2.632e-14
C119 1768 1803 2.871e-14
C117 1770 1803 6.85e-14
C115 1772 1803 2.321e-14
C114 1773 1803 4.869e-14
C113 1774 1803 5.165e-14
C112 1775 1803 7.43e-15
C111 1776 1803 2.455e-14
C109 1778 1803 6.107e-14
C108 1779 1803 2.785e-13
C107 1780 1803 4.11e-15
C104 1783 1803 1.96089e-12
C101 1786 1803 2.605e-14
C100 1787 1803 5.981e-14
C99 1788 1803 5.657e-14
C97 1790 1803 1.767e-14
C95 1792 1803 4.0891e-13
C93 1794 1803 2.596e-14
C90 1797 1803 5.1e-14
C89 1798 1803 1.662e-14
C88 1799 1803 1.198e-13
C86 1801 1803 2.16e-14
C84 1803 1803 2.08039e-11
C83 1804 1803 5.323e-14
C82 1805 1803 2.596e-14
C81 1806 1803 3.7515e-13
C80 1807 1803 9.7e-15
C79 1808 1803 2.16e-14
C78 1809 1803 4.881e-14
C77 1810 1803 1.8635e-14
C76 1811 1803 1.8635e-14
C75 1812 1803 4.678e-14
C74 1813 1803 5.578e-14
C73 1814 1803 4.768e-14
C72 1815 1803 2.299e-14
C70 1817 1803 8.58e-15
C69 1818 1803 4.686e-14
C67 1820 1803 5.521e-14
C65 1822 1803 2.871e-14
C64 1823 1803 2.005e-14
C63 1824 1803 8.53e-14
C61 1826 1803 2.321e-14
C59 1828 1803 2.632e-14
C58 1829 1803 5.165e-14
C57 1830 1803 4.869e-14
C56 1831 1803 3.2702e-13
C55 1832 1803 5.111e-14
C54 1833 1803 2.3943e-13
C52 1835 1803 1.8635e-14
C51 1836 1803 2.4045e-13
C50 1837 1803 3.9796e-13
C48 1839 1803 1.8635e-14
C47 1840 1803 4.66311e-13
C46 1841 1803 1.8635e-14
C45 1842 1803 4.8586e-13
C44 1843 1803 1.3724e-13
C42 1845 1803 2.74538e-12
C41 1846 1803 1.4596e-13
C40 1847 1803 1.8635e-14
C38 1849 1803 5.521e-14
C37 1850 1803 2.1294e-13
C36 1851 1803 1.8635e-14
C34 1853 1803 3.8105e-13
C33 1854 1803 1.8635e-14
C32 1855 1803 9.707e-14
C31 1856 1803 8.374e-14
C30 1857 1803 6.071e-14
C29 1858 1803 1.2737e-13
C26 1861 1803 3.7889e-13
C24 1863 1803 2.871e-14
C23 1864 1803 2.005e-14
C20 1867 1803 2.632e-14
C19 1868 1803 4.7371e-13
C18 1869 1803 6.378e-14
C17 1870 1803 2.321e-14
C16 1871 1803 5.165e-14
C15 1872 1803 4.869e-14
C14 1873 1803 5.38321e-13
C12 1875 1803 4.7044e-13
C11 1876 1803 2.871e-14
C10 1877 1803 2.005e-14
C8 1879 1803 2.632e-14
C7 1880 1803 7.206e-14
C6 1881 1803 2.87494e-12
C4 1883 1803 2.321e-14
C3 1884 1803 4.869e-14
C2 1885 1803 2.17515e-11
C1 1886 1803 5.165e-14
.ends act5_cougar

