* Spice description of mul2b_cougar
* Spice driver version -1209491804
* Date ( dd/mm/yyyy hh:mm:ss ):  9/10/2020 at 21:02:26

* INTERF vdd vss x[0] x[1] y[0] y[1] z[0] z[1] z[2] z[3] 


.subckt mul2b_cougar vdd vss x[0] x[1] y[0] y[1] z[0] z[1] z[2] z[3] 
Mtr_00188 sig13 rtl_map_3 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00187 vdd rtl_map_2 sig10 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00186 u0.y0.xr2_x1_sig sig13 sig11 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00185 sig11 rtl_map_2 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00184 sig11 sig10 u0.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00183 vdd rtl_map_3 sig11 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00182 cx[0] sig8 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00181 sig4 rtl_map_2 sig6 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00180 sig4 rtl_map_3 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00179 vdd rtl_map_2 sig4 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00178 sig6 rtl_map_3 sig8 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00177 sig8 u0.x1 sig4 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00176 sig17 u0.x1 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 vdd u0.y0.xr2_x1_sig sig14 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 sx[0] sig17 sig15 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00173 sig15 u0.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00172 sig15 sig14 sx[0] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00171 vdd u0.x1 sig15 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00170 z[0] sig19 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00169 vdd sx[0] sig19 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00168 sig27 u1.x1 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 vdd u1.y0.xr2_x1_sig sig22 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 sx[1] sig27 sig50 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00165 sig50 u1.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00164 sig50 sig22 sx[1] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00163 vdd u1.x1 sig50 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00162 sig31 rtl_map_1 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 vdd cx[0] sig29 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00160 u1.y0.xr2_x1_sig sig31 sig52 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00159 sig52 cx[0] vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00158 sig52 sig29 u1.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00157 vdd rtl_map_1 sig52 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00156 cx[1] sig37 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00155 sig53 cx[0] sig54 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00154 sig53 rtl_map_1 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00153 vdd cx[0] sig53 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00152 sig54 rtl_map_1 sig37 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00151 sig37 u1.x1 sig53 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00150 z[1] sig42 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00149 vdd sx[2] sig42 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00148 z[2] sig46 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00147 vdd sx[3] sig46 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00146 u1.x1 sig59 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00145 vdd y[0] sig59 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00144 sig59 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00143 u0.x1 sig60 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00142 vdd y[0] sig60 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 sig60 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 u3.x1 sig56 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00139 vdd y[1] sig56 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 sig56 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 cx[3] sig62 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00136 sig64 cx[2] sig63 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00135 sig64 cx[1] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00134 vdd cx[2] sig64 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00133 sig63 cx[1] sig62 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00132 sig62 u3.x1 sig64 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00131 sig69 cx[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00130 vdd cx[2] sig66 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 u3.y0.xr2_x1_sig sig69 sig67 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00128 sig67 cx[2] vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00127 sig67 sig66 u3.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00126 vdd cx[1] sig67 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00125 sig72 u3.x1 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 vdd u3.y0.xr2_x1_sig sig71 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00123 sx[3] sig72 sig70 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00122 sig70 u3.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00121 sig70 sig71 sx[3] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00120 vdd u3.x1 sig70 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00119 u2.x1 sig77 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00118 vdd y[1] sig77 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 sig77 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 sig88 sx[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 vdd rtl_map_0 sig87 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 u2.y0.xr2_x1_sig sig88 sig104 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00113 sig104 rtl_map_0 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00112 sig104 sig87 u2.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00111 vdd sx[1] sig104 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00110 sig94 u2.x1 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 vdd u2.y0.xr2_x1_sig sig93 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 sx[2] sig94 sig105 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00107 sig105 u2.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00106 sig105 sig93 sx[2] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00105 vdd u2.x1 sig105 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00104 z[3] sig98 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00103 vdd cx[3] sig98 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00102 cx[2] sig80 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00101 sig102 rtl_map_0 sig103 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00100 sig102 sx[1] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00099 vdd rtl_map_0 sig102 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00098 sig103 sx[1] sig80 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00097 sig80 u2.x1 sig102 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00096 vss vdd rtl_map_3 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00095 sig10 rtl_map_2 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00094 vss rtl_map_3 sig13 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00093 sig38 sig13 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00092 u0.y0.xr2_x1_sig sig10 sig38 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 sig35 rtl_map_3 u0.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 vss rtl_map_2 sig35 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 vss sig8 cx[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 vss rtl_map_3 sig30 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00087 sig30 rtl_map_2 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00086 sig8 rtl_map_3 sig28 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00085 sig28 rtl_map_2 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00084 sig30 u0.x1 sig8 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00083 sig14 u0.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00082 vss u0.x1 sig17 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00081 sig44 sig17 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 sx[0] sig14 sig44 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 sig41 u0.x1 sx[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 vss u0.y0.xr2_x1_sig sig41 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 vss vdd rtl_map_2 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00076 vss sig19 z[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00075 sig19 sx[0] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00074 sig22 u1.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00073 vss u1.x1 sig27 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00072 sig21 sig27 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 sx[1] sig22 sig21 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 sig23 u1.x1 sx[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 vss u1.y0.xr2_x1_sig sig23 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 sig29 cx[0] vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00067 vss rtl_map_1 sig31 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00066 sig33 sig31 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 u1.y0.xr2_x1_sig sig29 sig33 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 sig32 rtl_map_1 u1.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 vss cx[0] sig32 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 vss sig37 cx[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 vss rtl_map_1 sig39 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00060 sig39 cx[0] vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00059 sig37 rtl_map_1 sig36 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00058 sig36 cx[0] vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00057 sig39 u1.x1 sig37 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00056 vss sig42 z[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 sig42 sx[2] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00054 vss sig46 z[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 sig46 sx[3] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00052 vss vdd rtl_map_1 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00051 sig59 x[1] sig78 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 vss sig59 u1.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 sig78 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 sig60 x[0] sig79 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 vss sig60 u0.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 sig79 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 sig56 x[1] sig73 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 vss sig56 u3.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 sig73 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 vss sig62 cx[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 vss cx[1] sig81 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00040 sig81 cx[2] vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00039 sig62 cx[1] sig82 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00038 sig82 cx[2] vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00037 sig81 u3.x1 sig62 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00036 sig66 cx[2] vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00035 vss cx[1] sig69 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 sig89 sig69 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 u3.y0.xr2_x1_sig sig66 sig89 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 sig91 cx[1] u3.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 vss cx[2] sig91 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 sig71 u3.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 vss u3.x1 sig72 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 sig95 sig72 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 sx[3] sig71 sig95 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 sig96 u3.x1 sx[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 vss u3.y0.xr2_x1_sig sig96 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 sig77 x[0] sig76 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 vss sig77 u2.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 sig76 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 sig87 rtl_map_0 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 vss sx[1] sig88 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00019 sig85 sig88 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 u2.y0.xr2_x1_sig sig87 sig85 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 sig83 sx[1] u2.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 vss rtl_map_0 sig83 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 sig93 u2.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 vss u2.x1 sig94 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 sig90 sig94 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 sx[2] sig93 sig90 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 sig92 u2.x1 sx[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 vss u2.y0.xr2_x1_sig sig92 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 vss sig98 z[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 sig98 cx[3] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00007 vss vdd rtl_map_0 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 vss sig80 cx[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 vss sx[1] sig100 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00004 sig100 rtl_map_0 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00003 sig80 sx[1] sig101 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00002 sig101 rtl_map_0 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00001 sig100 u2.x1 sig80 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
C105 sig105 vss 9.7e-15
C104 sig104 vss 9.7e-15
C102 sig102 vss 8.58e-15
C100 sig100 vss 4.11e-15
C98 sig98 vss 1.568e-14
C97 z[3] vss 2.659e-14
C94 sig94 vss 2.596e-14
C93 sig93 vss 2.16e-14
C88 sig88 vss 2.596e-14
C87 sig87 vss 2.16e-14
C86 rtl_map_0 vss 1.0243e-13
C84 u2.y0.xr2_x1_sig vss 5.991e-14
C81 sig81 vss 4.11e-15
C80 sig80 vss 2.299e-14
C77 sig77 vss 1.8635e-14
C75 u2.x1 vss 1.0949e-13
C72 sig72 vss 2.596e-14
C71 sig71 vss 2.16e-14
C70 sig70 vss 9.7e-15
C69 sig69 vss 2.596e-14
C68 u3.y0.xr2_x1_sig vss 5.751e-14
C67 sig67 vss 9.7e-15
C66 sig66 vss 2.16e-14
C65 cx[3] vss 7.301e-14
C64 sig64 vss 8.58e-15
C62 sig62 vss 2.299e-14
C61 cx[2] vss 1.1155e-13
C60 sig60 vss 1.8635e-14
C59 sig59 vss 1.8635e-14
C58 y[0] vss 8.493e-14
C57 y[1] vss 7.197e-14
C56 sig56 vss 1.8635e-14
C55 u3.x1 vss 1.1909e-13
C53 sig53 vss 8.58e-15
C52 sig52 vss 9.7e-15
C51 x[1] vss 5.257e-14
C50 sig50 vss 9.7e-15
C49 sx[3] vss 5.859e-14
C48 z[2] vss 3.427e-14
C47 sx[2] vss 7.179e-14
C46 sig46 vss 1.568e-14
C45 z[1] vss 3.259e-14
C42 sig42 vss 1.568e-14
C40 cx[1] vss 1.1768e-13
C39 sig39 vss 4.11e-15
C37 sig37 vss 2.299e-14
C34 rtl_map_1 vss 1.0392e-13
C31 sig31 vss 2.596e-14
C30 sig30 vss 4.11e-15
C29 sig29 vss 2.16e-14
C27 sig27 vss 2.596e-14
C26 u1.x1 vss 1.0301e-13
C25 u1.y0.xr2_x1_sig vss 6.351e-14
C24 sx[1] vss 1.371e-13
C22 sig22 vss 2.16e-14
C20 vss vss 1.1514e-12
C19 sig19 vss 1.568e-14
C18 z[0] vss 2.371e-14
C17 sig17 vss 2.596e-14
C16 sx[0] vss 5.859e-14
C15 sig15 vss 9.7e-15
C14 sig14 vss 2.16e-14
C13 sig13 vss 2.596e-14
C12 u0.y0.xr2_x1_sig vss 5.991e-14
C11 sig11 vss 9.7e-15
C10 sig10 vss 2.16e-14
C9 u0.x1 vss 1.2269e-13
C8 sig8 vss 2.299e-14
C7 cx[0] vss 1.2147e-13
C5 rtl_map_2 vss 1.0603e-13
C4 sig4 vss 8.58e-15
C3 x[0] vss 9.481e-14
C2 rtl_map_3 vss 1.1472e-13
C1 vdd vss 1.22168e-12
.ends mul2b_cougar

