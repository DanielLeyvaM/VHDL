* Spice description of sum3b_cougar
* Spice driver version -1208947036
* Date ( dd/mm/yyyy hh:mm:ss ): 26/10/2020 at 21:03:50

* INTERF a[0] a[1] a[2] b[0] b[1] b[2] ci co so[0] so[1] so[2] vdd vss 


.subckt sum3b_cougar 62 42 18 61 56 54 57 14 52 30 9 66 49 
* NET 9 = so[2]
* NET 14 = co
* NET 18 = a[2]
* NET 20 = xr2_x1_3_sig
* NET 28 = mbk_buf_aux4
* NET 30 = so[1]
* NET 35 = aux7
* NET 36 = a2_x2_sig
* NET 42 = a[1]
* NET 43 = xr2_x1_2_sig
* NET 49 = vss
* NET 52 = so[0]
* NET 54 = b[2]
* NET 55 = aux4
* NET 56 = b[1]
* NET 57 = ci
* NET 61 = b[0]
* NET 62 = a[0]
* NET 65 = xr2_x1_sig
* NET 66 = vdd
Mtr_00116 55 58 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00115 60 61 59 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00114 60 62 66 66 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00113 66 61 60 66 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00112 59 62 58 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00111 58 57 60 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00110 63 62 66 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 66 61 64 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 65 63 67 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00107 67 61 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00106 67 64 65 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00105 66 62 67 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00104 50 57 66 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 66 65 51 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 52 50 53 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00101 53 65 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00100 53 51 52 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00099 66 57 53 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00098 41 56 66 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 66 42 45 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 43 41 26 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00095 26 42 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00094 26 45 43 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00093 66 56 26 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00092 25 55 66 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 24 42 38 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 66 56 24 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 38 36 25 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 35 38 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00087 27 43 66 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 66 28 33 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 30 27 23 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00084 23 28 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00083 23 33 30 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00082 66 43 23 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00081 19 18 66 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 66 54 22 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 20 19 21 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00078 21 54 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00077 21 22 20 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00076 66 18 21 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00075 14 16 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00074 15 54 12 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00073 15 18 66 66 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00072 66 54 15 66 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00071 12 18 16 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00070 16 35 15 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00069 8 20 66 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 66 35 10 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 9 8 11 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00066 11 35 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00065 11 10 9 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00064 66 20 11 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00063 28 13 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00062 66 55 13 66 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00061 36 17 66 66 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00060 66 42 17 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 17 56 66 66 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 49 58 55 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 49 62 40 49 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00056 40 61 49 49 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00055 58 62 39 49 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00054 39 61 49 49 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00053 40 57 58 49 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00052 64 61 49 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00051 49 62 63 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00050 47 63 49 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 65 64 47 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 48 62 65 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 49 61 48 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 51 65 49 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 49 57 50 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00044 34 50 49 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 52 51 34 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 32 57 52 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 49 65 32 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 45 42 49 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00039 49 56 41 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 46 41 49 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 43 45 46 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 44 56 43 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 49 42 44 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 37 42 49 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 49 56 37 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 37 55 38 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00031 38 36 37 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00030 49 38 35 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 33 28 49 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 49 43 27 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00027 29 27 49 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 30 33 29 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 31 43 30 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 49 28 31 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 22 54 49 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 49 18 19 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00021 7 19 49 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 20 22 7 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 6 18 20 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 49 54 6 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 49 16 14 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 49 18 4 49 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00015 4 54 49 49 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00014 16 18 3 49 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00013 3 54 49 49 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00012 4 35 16 49 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00011 10 35 49 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 49 20 8 49 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 1 8 49 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 9 10 1 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 2 20 9 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 49 35 2 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 49 13 28 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 13 55 49 49 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00003 17 56 5 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 49 17 36 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 5 42 49 49 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C66 4 49 4.11e-15
C61 8 49 2.596e-14
C60 9 49 3.409e-14
C59 10 49 2.16e-14
C58 11 49 9.7e-15
C56 13 49 1.568e-14
C55 14 49 3.344e-14
C54 15 49 8.58e-15
C53 16 49 2.299e-14
C52 17 49 1.8635e-14
C51 18 49 8.803e-14
C50 19 49 2.596e-14
C49 20 49 9.115e-14
C48 21 49 9.7e-15
C47 22 49 2.16e-14
C46 23 49 9.7e-15
C42 26 49 9.7e-15
C41 27 49 2.596e-14
C40 28 49 5.649e-14
C38 30 49 3.649e-14
C35 33 49 2.16e-14
C33 35 49 9.793e-14
C32 36 49 5.143e-14
C31 37 49 7.43e-15
C30 38 49 2.639e-14
C28 40 49 4.11e-15
C27 41 49 2.596e-14
C26 42 49 1.086e-13
C25 43 49 8.995e-14
C23 45 49 2.16e-14
C19 49 49 6.42961e-13
C18 50 49 2.596e-14
C17 51 49 2.16e-14
C16 52 49 3.649e-14
C15 53 49 9.7e-15
C14 54 49 1.2851e-13
C13 55 49 1.0326e-13
C12 56 49 1.2001e-13
C11 57 49 1.1309e-13
C10 58 49 2.299e-14
C8 60 49 8.58e-15
C7 61 49 9.979e-14
C6 62 49 9.531e-14
C5 63 49 2.596e-14
C4 64 49 2.16e-14
C3 65 49 8.271e-14
C2 66 49 6.55001e-13
C1 67 49 9.7e-15
.ends sum3b_cougar

