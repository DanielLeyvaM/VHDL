* Spice description of mul5b_cougar
* Spice driver version -1209295196
* Date ( dd/mm/yyyy hh:mm:ss ):  4/11/2020 at 11:15:31

* INTERF vdd vss x[0] x[1] x[2] x[3] x[4] y[0] y[1] y[2] y[3] y[4] z[0] z[1] 
* INTERF z[2] z[3] z[4] z[5] z[6] z[7] z[8] z[9] 


.subckt mul5b_cougar vdd vss x[0] x[1] x[2] x[3] x[4] y[0] y[1] y[2] y[3] y[4] z[0] z[1] z[2] z[3] z[4] z[5] z[6] z[7] z[8] z[9] 
Mtr_01100 u5.x1 sig3 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01099 vdd y[1] sig3 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01098 sig3 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01097 cx[5] sig15 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01096 sig12 u5.x1 sig13 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01095 sig12 rtl_map_3 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01094 vdd u5.x1 sig12 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01093 sig13 rtl_map_3 sig15 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01092 sig15 sx[1] sig12 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01091 sig9 rtl_map_3 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01090 vdd u5.x1 sig8 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01089 u5.y0.xr2_x1_sig sig9 sig10 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01088 sig10 u5.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01087 sig10 sig8 u5.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01086 vdd rtl_map_3 sig10 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01085 sig29 rtl_map_2 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01084 vdd u10.x1 sig26 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01083 u10.y0.xr2_x1_sig sig29 sig27 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01082 sig27 u10.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01081 sig27 sig26 u10.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01080 vdd rtl_map_2 sig27 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01079 u10.x1 sig17 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01078 vdd y[2] sig17 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01077 sig17 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01076 cx[10] sig22 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01075 sig19 u10.x1 sig21 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01074 sig19 rtl_map_2 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01073 vdd u10.x1 sig19 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01072 sig21 rtl_map_2 sig22 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01071 sig22 sx[6] sig19 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01070 sig33 sx[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01069 vdd u5.y0.xr2_x1_sig sig32 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01068 sx[5] sig33 sig30 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01067 sig30 u5.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01066 sig30 sig32 sx[5] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01065 vdd sx[1] sig30 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01064 z[0] sig37 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01063 vdd sx[0] sig37 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01062 z[1] sig35 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01061 vdd sx[5] sig35 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01060 sig50 cx[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01059 vdd u3.x1 sig47 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01058 u3.y0.xr2_x1_sig sig50 sig100 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01057 sig100 u3.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01056 sig100 sig47 u3.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01055 vdd cx[2] sig100 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01054 sig45 rtl_map_5 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01053 vdd u3.y0.xr2_x1_sig sig40 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01052 sx[3] sig45 sig99 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01051 sig99 u3.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01050 sig99 sig40 sx[3] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01049 vdd rtl_map_5 sig99 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01048 cx[6] sig57 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01047 sig101 u6.x1 sig102 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01046 sig101 cx[5] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01045 vdd u6.x1 sig101 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01044 sig102 cx[5] sig57 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01043 sig57 sx[2] sig101 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01042 sig64 cx[5] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01041 vdd u6.x1 sig61 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01040 u6.y0.xr2_x1_sig sig64 sig103 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01039 sig103 u6.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01038 sig103 sig61 u6.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01037 vdd cx[5] sig103 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01036 sig86 sx[6] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01035 vdd u10.y0.xr2_x1_sig sig84 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01034 sx[10] sig86 sig106 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01033 sig106 u10.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01032 sig106 sig84 sx[10] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01031 vdd sx[6] sig106 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01030 sig71 sx[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01029 vdd u6.y0.xr2_x1_sig sig69 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01028 sx[6] sig71 sig104 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01027 sig104 u6.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01026 sig104 sig69 sx[6] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01025 vdd sx[2] sig104 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01024 sig81 rtl_map_7 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01023 vdd u1.y0.xr2_x1_sig sig78 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01022 sx[1] sig81 sig105 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01021 sig105 u1.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01020 sig105 sig78 sx[1] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01019 vdd rtl_map_7 sig105 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01018 z[2] sig90 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01017 vdd sx[10] sig90 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01016 sig98 rtl_map_9 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01015 vdd u0.y0.xr2_x1_sig sig95 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01014 sx[0] sig98 sig107 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01013 sig107 u0.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01012 sig107 sig95 sx[0] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01011 vdd rtl_map_9 sig107 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01010 cx[3] sig110 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01009 sig108 u3.x1 sig109 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01008 sig108 cx[2] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01007 vdd u3.x1 sig108 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01006 sig109 cx[2] sig110 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01005 sig110 rtl_map_5 sig108 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01004 u3.x1 sig112 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01003 vdd y[0] sig112 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01002 sig112 x[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01001 cx[2] sig119 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01000 sig115 u2.x1 sig118 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00999 sig115 cx[1] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00998 vdd u2.x1 sig115 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00997 sig118 cx[1] sig119 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00996 sig119 rtl_map_6 sig115 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00995 sig127 cx[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00994 vdd u2.x1 sig125 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00993 u2.y0.xr2_x1_sig sig127 sig126 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00992 sig126 u2.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00991 sig126 sig125 u2.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00990 vdd cx[1] sig126 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00989 sig123 rtl_map_6 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00988 vdd u2.y0.xr2_x1_sig sig121 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00987 sx[2] sig123 sig124 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00986 sig124 u2.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00985 sig124 sig121 sx[2] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00984 vdd rtl_map_6 sig124 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00983 cx[1] sig128 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00982 sig129 u1.x1 sig132 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00981 sig129 cx[0] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00980 vdd u1.x1 sig129 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00979 sig132 cx[0] sig128 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00978 sig128 rtl_map_7 sig129 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00977 u0.x1 sig137 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00976 vdd y[0] sig137 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00975 sig137 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00974 sig135 cx[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00973 vdd u1.x1 sig134 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00972 u1.y0.xr2_x1_sig sig135 sig133 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00971 sig133 u1.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00970 sig133 sig134 u1.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00969 vdd cx[0] sig133 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00968 sig144 rtl_map_8 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00967 vdd u0.x1 sig143 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00966 u0.y0.xr2_x1_sig sig144 sig142 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00965 sig142 u0.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00964 sig142 sig143 u0.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00963 vdd rtl_map_8 sig142 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00962 cx[0] sig140 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00961 sig138 u0.x1 sig139 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00960 sig138 rtl_map_8 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00959 vdd u0.x1 sig138 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00958 sig139 rtl_map_8 sig140 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00957 sig140 rtl_map_9 sig138 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00956 sig156 cx[6] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00955 vdd u7.x1 sig155 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00954 u7.y0.xr2_x1_sig sig156 sig216 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00953 sig216 u7.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00952 sig216 sig155 u7.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00951 vdd cx[6] sig216 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00950 sig162 sx[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00949 vdd u7.y0.xr2_x1_sig sig163 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00948 sx[7] sig162 sig217 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00947 sig217 u7.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00946 sig217 sig163 sx[7] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00945 vdd sx[3] sig217 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00944 cx[7] sig149 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00943 sig212 u7.x1 sig214 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00942 sig212 cx[6] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00941 vdd u7.x1 sig212 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00940 sig214 cx[6] sig149 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00939 sig149 sx[3] sig212 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00938 u2.x1 sig169 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00937 vdd y[0] sig169 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00936 sig169 x[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00935 u16.x1 sig175 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00934 vdd y[3] sig175 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00933 sig175 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00932 u15.x1 sig183 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00931 vdd y[3] sig183 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00930 sig183 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00929 u6.x1 sig165 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00928 vdd y[1] sig165 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00927 sig165 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00926 sig190 rtl_map_1 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00925 vdd u15.x1 sig192 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00924 u15.y0.xr2_x1_sig sig190 sig223 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00923 sig223 u15.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00922 sig223 sig192 u15.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00921 vdd rtl_map_1 sig223 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00920 cx[15] sig184 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00919 sig219 u15.x1 sig221 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00918 sig219 rtl_map_1 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00917 vdd u15.x1 sig219 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00916 sig221 rtl_map_1 sig184 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00915 sig184 sx[11] sig219 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00914 u20.x1 sig197 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00913 vdd y[4] sig197 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00912 sig197 x[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00911 sig206 sx[11] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00910 vdd u15.y0.xr2_x1_sig sig205 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00909 sx[15] sig206 sig225 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00908 sig225 u15.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00907 sig225 sig205 sx[15] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00906 vdd sx[11] sig225 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00905 u1.x1 sig178 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00904 vdd y[0] sig178 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00903 sig178 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00902 z[3] sig209 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00901 vdd sx[15] sig209 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00900 u7.x1 sig232 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00899 vdd y[1] sig232 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00898 sig232 x[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00897 u8.x1 sig226 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00896 vdd y[1] sig226 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00895 sig226 x[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00894 sig231 cx[7] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00893 vdd u8.x1 sig228 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00892 u8.y0.xr2_x1_sig sig231 sig230 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00891 sig230 u8.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00890 sig230 sig228 u8.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00889 vdd cx[7] sig230 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00888 sig243 cx[15] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00887 vdd u16.x1 sig242 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00886 u16.y0.xr2_x1_sig sig243 sig241 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00885 sig241 u16.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00884 sig241 sig242 u16.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00883 vdd cx[15] sig241 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00882 cx[16] sig237 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00881 sig235 u16.x1 sig236 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00880 sig235 cx[15] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00879 vdd u16.x1 sig235 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00878 sig236 cx[15] sig237 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00877 sig237 sx[12] sig235 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00876 u11.x1 sig233 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00875 vdd y[2] sig233 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00874 sig233 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00873 sig245 sx[12] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00872 vdd u16.y0.xr2_x1_sig sig244 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00871 sx[16] sig245 sig246 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00870 sig246 u16.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00869 sig246 sig244 sx[16] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00868 vdd sx[12] sig246 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00867 u21.x1 sig248 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00866 vdd y[4] sig248 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00865 sig248 x[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00864 cx[20] sig252 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00863 sig249 u20.x1 sig253 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00862 sig249 rtl_map_0 vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00861 vdd u20.x1 sig249 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00860 sig253 rtl_map_0 sig252 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00859 sig252 sx[16] sig249 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00858 sig257 rtl_map_0 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00857 vdd u20.x1 sig255 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00856 u20.y0.xr2_x1_sig sig257 sig254 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00855 sig254 u20.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00854 sig254 sig255 u20.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00853 vdd rtl_map_0 sig254 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00852 sig261 sx[16] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00851 vdd u20.y0.xr2_x1_sig sig258 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00850 sx[20] sig261 sig260 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00849 sig260 u20.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00848 sig260 sig258 sx[20] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00847 vdd sx[16] sig260 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00846 z[4] sig262 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00845 vdd sx[20] sig262 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00844 cx[8] sig306 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00843 sig310 u8.x1 sig311 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00842 sig310 cx[7] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00841 vdd u8.x1 sig310 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00840 sig311 cx[7] sig306 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00839 sig306 sx[4] sig310 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00838 sig269 sx[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00837 vdd u8.y0.xr2_x1_sig sig268 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00836 sx[8] sig269 sig315 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00835 sig315 u8.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00834 sig315 sig268 sx[8] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00833 vdd sx[4] sig315 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00832 sig273 cx[11] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00831 vdd u12.x1 sig276 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00830 u12.y0.xr2_x1_sig sig273 sig318 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00829 sig318 u12.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00828 sig318 sig276 u12.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00827 vdd cx[11] sig318 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00826 sig282 sx[8] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00825 vdd u12.y0.xr2_x1_sig sig281 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00824 sx[12] sig282 sig320 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00823 sig320 u12.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00822 sig320 sig281 sx[12] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00821 vdd sx[8] sig320 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00820 sig288 cx[10] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00819 vdd u11.x1 sig287 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00818 u11.y0.xr2_x1_sig sig288 sig329 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00817 sig329 u11.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00816 sig329 sig287 u11.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00815 vdd cx[10] sig329 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00814 cx[11] sig322 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00813 sig325 u11.x1 sig326 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00812 sig325 cx[10] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00811 vdd u11.x1 sig325 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00810 sig326 cx[10] sig322 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00809 sig322 sx[7] sig325 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00808 sig293 sx[7] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00807 vdd u11.y0.xr2_x1_sig sig292 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00806 sx[11] sig293 sig331 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00805 sig331 u11.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00804 sig331 sig292 sx[11] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00803 vdd sx[7] sig331 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00802 sig298 cx[20] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00801 vdd u21.x1 sig297 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00800 u21.y0.xr2_x1_sig sig298 sig340 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00799 sig340 u21.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00798 sig340 sig297 u21.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00797 vdd cx[20] sig340 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00796 cx[21] sig334 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00795 sig333 u21.x1 sig337 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00794 sig333 cx[20] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00793 vdd u21.x1 sig333 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00792 sig337 cx[20] sig334 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00791 sig334 sx[17] sig333 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00790 sig302 sx[17] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00789 vdd u21.y0.xr2_x1_sig sig301 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00788 sx[21] sig302 sig345 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00787 sig345 u21.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00786 sig345 sig301 sx[21] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00785 vdd sx[17] sig345 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00784 z[5] sig305 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00783 vdd sx[21] sig305 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00782 sig351 rtl_map_4 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00781 vdd u4.y0.xr2_x1_sig sig348 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00780 sx[4] sig351 sig347 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00779 sig347 u4.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00778 sig347 sig348 sx[4] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00777 vdd rtl_map_4 sig347 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00776 u12.x1 sig352 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00775 vdd y[2] sig352 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00774 sig352 x[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00773 cx[12] sig356 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00772 sig353 u12.x1 sig354 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00771 sig353 cx[11] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00770 vdd u12.x1 sig353 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00769 sig354 cx[11] sig356 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00768 sig356 sx[8] sig353 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00767 u17.x1 sig357 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00766 vdd y[3] sig357 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00765 sig357 x[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00764 sig370 sx[13] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00763 vdd u17.y0.xr2_x1_sig sig369 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00762 sx[17] sig370 sig368 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00761 sig368 u17.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00760 sig368 sig369 sx[17] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00759 vdd sx[13] sig368 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00758 sig367 cx[16] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00757 vdd u17.x1 sig364 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00756 u17.y0.xr2_x1_sig sig367 sig363 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00755 sig363 u17.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00754 sig363 sig364 u17.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00753 vdd cx[16] sig363 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00752 cx[17] sig361 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00751 sig359 u17.x1 sig360 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00750 sig359 cx[16] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00749 vdd u17.x1 sig359 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00748 sig360 cx[16] sig361 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00747 sig361 sx[13] sig359 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00746 u22.x1 sig371 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00745 vdd y[4] sig371 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00744 sig371 x[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00743 sig376 cx[21] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00742 vdd u22.x1 sig374 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00741 u22.y0.xr2_x1_sig sig376 sig373 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00740 sig373 u22.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00739 sig373 sig374 u22.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00738 vdd cx[21] sig373 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00737 z[6] sig383 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00736 vdd sx[22] sig383 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00735 sig381 sx[18] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00734 vdd u22.y0.xr2_x1_sig sig377 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00733 sx[22] sig381 sig378 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00732 sig378 u22.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00731 sig378 sig377 sx[22] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00730 vdd sx[18] sig378 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00729 sig405 cx[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00728 vdd u4.x1 sig402 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00727 u4.y0.xr2_x1_sig sig405 sig449 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00726 sig449 u4.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00725 sig449 sig402 u4.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00724 vdd cx[3] sig449 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00723 cx[4] sig408 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00722 sig456 u4.x1 sig458 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00721 sig456 cx[3] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00720 vdd u4.x1 sig456 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00719 sig458 cx[3] sig408 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00718 sig408 rtl_map_4 sig456 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00717 sig421 sx[9] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00716 vdd u13.y0.xr2_x1_sig sig420 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00715 sx[13] sig421 sig468 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00714 sig468 u13.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00713 sig468 sig420 sx[13] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00712 vdd sx[9] sig468 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00711 u13.x1 sig410 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00710 vdd y[2] sig410 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00709 sig410 x[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00708 sig415 cx[12] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00707 vdd u13.x1 sig414 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00706 u13.y0.xr2_x1_sig sig415 sig465 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00705 sig465 u13.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00704 sig465 sig414 u13.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00703 vdd cx[12] sig465 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00702 sig435 cx[17] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00701 vdd u18.x1 sig434 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00700 u18.y0.xr2_x1_sig sig435 sig485 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00699 sig485 u18.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00698 sig485 sig434 u18.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00697 vdd cx[17] sig485 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00696 u18.x1 sig430 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00695 vdd y[3] sig430 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00694 sig430 x[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00693 cx[18] sig424 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00692 sig475 u18.x1 sig481 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00691 sig475 cx[17] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00690 vdd u18.x1 sig475 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00689 sig481 cx[17] sig424 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00688 sig424 sx[14] sig475 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00687 sig442 sx[14] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00686 vdd u18.y0.xr2_x1_sig sig440 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00685 sx[18] sig442 sig500 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00684 sig500 u18.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00683 sig500 sig440 sx[18] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00682 vdd sx[14] sig500 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00681 cx[22] sig437 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00680 sig491 u22.x1 sig492 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00679 sig491 cx[21] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00678 vdd u22.x1 sig491 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00677 sig492 cx[21] sig437 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00676 sig437 sx[18] sig491 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00675 z[7] sig446 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00674 vdd sx[23] sig446 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00673 u4.x1 sig455 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00672 vdd y[0] sig455 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00671 sig455 x[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00670 sig454 cx[8] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00669 vdd u9.x1 sig451 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00668 u9.y0.xr2_x1_sig sig454 sig450 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00667 sig450 u9.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00666 sig450 sig451 u9.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00665 vdd cx[8] sig450 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00664 sig461 cx[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00663 vdd u9.y0.xr2_x1_sig sig459 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00662 sx[9] sig461 sig460 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00661 sig460 u9.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00660 sig460 sig459 sx[9] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00659 vdd cx[4] sig460 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00658 u19.x1 sig466 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00657 vdd y[3] sig466 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00656 sig466 x[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00655 cx[13] sig463 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00654 sig464 u13.x1 sig462 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00653 sig464 cx[12] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00652 vdd u13.x1 sig464 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00651 sig462 cx[12] sig463 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00650 sig463 sx[9] sig464 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00649 cx[19] sig472 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00648 sig470 u19.x1 sig473 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00647 sig470 cx[18] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00646 vdd u19.x1 sig470 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00645 sig473 cx[18] sig472 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00644 sig472 cx[14] sig470 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00643 sig483 cx[14] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00642 vdd u19.y0.xr2_x1_sig sig480 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00641 sx[19] sig483 sig482 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00640 sig482 u19.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00639 sig482 sig480 sx[19] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00638 vdd cx[14] sig482 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00637 sig479 cx[18] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00636 vdd u19.x1 sig478 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00635 u19.y0.xr2_x1_sig sig479 sig476 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00634 sig476 u19.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00633 sig476 sig478 u19.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00632 vdd cx[18] sig476 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00631 u24.x1 sig487 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00630 vdd y[4] sig487 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00629 sig487 x[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00628 u23.x1 sig488 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00627 vdd y[4] sig488 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00626 sig488 x[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00625 sig499 cx[22] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00624 vdd u23.x1 sig497 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00623 u23.y0.xr2_x1_sig sig499 sig496 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00622 sig496 u23.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00621 sig496 sig497 u23.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00620 vdd cx[22] sig496 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00619 cx[23] sig495 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00618 sig490 u23.x1 sig493 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00617 sig490 cx[22] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00616 vdd u23.x1 sig490 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00615 sig493 cx[22] sig495 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00614 sig495 sx[19] sig490 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00613 sig503 sx[19] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00612 vdd u23.y0.xr2_x1_sig sig501 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00611 sx[23] sig503 sig502 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00610 sig502 u23.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00609 sig502 sig501 sx[23] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00608 vdd sx[19] sig502 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00607 cx[9] sig530 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00606 sig568 u9.x1 sig567 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00605 sig568 cx[8] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00604 vdd u9.x1 sig568 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00603 sig567 cx[8] sig530 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00602 sig530 cx[4] sig568 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00601 u9.x1 sig528 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00600 vdd y[1] sig528 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00599 sig528 x[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00598 u14.x1 sig536 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00597 vdd y[2] sig536 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00596 sig536 x[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00595 sig544 cx[13] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00594 vdd u14.x1 sig540 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00593 u14.y0.xr2_x1_sig sig544 sig571 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00592 sig571 u14.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00591 sig571 sig540 u14.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00590 vdd cx[13] sig571 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00589 sig548 cx[9] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00588 vdd u14.y0.xr2_x1_sig sig546 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00587 sx[14] sig548 sig572 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00586 sig572 u14.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00585 sig572 sig546 sx[14] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00584 vdd cx[9] sig572 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00583 cx[14] sig537 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00582 sig569 u14.x1 sig570 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00581 sig569 cx[13] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00580 vdd u14.x1 sig569 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00579 sig570 cx[13] sig537 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00578 sig537 cx[9] sig569 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00577 cx[24] sig560 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00576 sig576 u24.x1 sig575 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00575 sig576 cx[23] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00574 vdd u24.x1 sig576 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00573 sig575 cx[23] sig560 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00572 sig560 cx[19] sig576 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00571 sig557 cx[23] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00570 vdd u24.x1 sig556 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00569 u24.y0.xr2_x1_sig sig557 sig574 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00568 sig574 u24.x1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00567 sig574 sig556 u24.y0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00566 vdd cx[23] sig574 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00565 z[8] sig563 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00564 vdd sx[24] sig563 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00563 z[9] sig565 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00562 vdd cx[24] sig565 vdd tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00561 sig552 cx[19] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00560 vdd u24.y0.xr2_x1_sig sig549 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00559 sx[24] sig552 sig573 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00558 sig573 u24.y0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00557 sig573 sig549 sx[24] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00556 vdd cx[19] sig573 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00555 sig3 x[0] sig46 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00554 vss sig3 u5.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00553 sig46 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00552 vss vdd rtl_map_5 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00551 vss vdd rtl_map_3 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00550 vss sig15 cx[5] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00549 vss rtl_map_3 sig63 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00548 sig63 u5.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00547 sig15 rtl_map_3 sig60 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00546 sig60 u5.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00545 sig63 sx[1] sig15 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00544 sig8 u5.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00543 vss rtl_map_3 sig9 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00542 sig54 sig9 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00541 u5.y0.xr2_x1_sig sig8 sig54 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00540 sig55 rtl_map_3 u5.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00539 vss u5.x1 sig55 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00538 sig26 u10.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00537 vss rtl_map_2 sig29 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00536 sig82 sig29 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00535 u10.y0.xr2_x1_sig sig26 sig82 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00534 sig83 rtl_map_2 u10.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00533 vss u10.x1 sig83 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00532 sig17 x[0] sig70 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00531 vss sig17 u10.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00530 sig70 y[2] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00529 vss sig22 cx[10] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00528 vss rtl_map_2 sig73 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00527 sig73 u10.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00526 sig22 rtl_map_2 sig74 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00525 sig74 u10.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00524 sig73 sx[6] sig22 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00523 vss vdd rtl_map_2 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00522 sig32 u5.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00521 vss sx[1] sig33 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00520 sig92 sig33 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00519 sx[5] sig32 sig92 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00518 sig89 sx[1] sx[5] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00517 vss u5.y0.xr2_x1_sig sig89 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00516 vss sig37 z[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00515 sig37 sx[0] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00514 vss sig35 z[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00513 sig35 sx[5] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00512 sig47 u3.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00511 vss cx[2] sig50 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00510 sig49 sig50 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00509 u3.y0.xr2_x1_sig sig47 sig49 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00508 sig51 cx[2] u3.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00507 vss u3.x1 sig51 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00506 sig40 u3.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00505 vss rtl_map_5 sig45 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00504 sig43 sig45 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00503 sx[3] sig40 sig43 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00502 sig41 rtl_map_5 sx[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00501 vss u3.y0.xr2_x1_sig sig41 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00500 vss sig57 cx[6] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00499 vss cx[5] sig56 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00498 sig56 u6.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00497 sig57 cx[5] sig58 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00496 sig58 u6.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00495 sig56 sx[2] sig57 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00494 sig61 u6.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00493 vss cx[5] sig64 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00492 sig67 sig64 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00491 u6.y0.xr2_x1_sig sig61 sig67 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00490 sig65 cx[5] u6.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00489 vss u6.x1 sig65 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00488 sig84 u10.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00487 vss sx[6] sig86 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00486 sig85 sig86 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00485 sx[10] sig84 sig85 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00484 sig87 sx[6] sx[10] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00483 vss u10.y0.xr2_x1_sig sig87 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00482 sig69 u6.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00481 vss sx[2] sig71 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00480 sig72 sig71 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00479 sx[6] sig69 sig72 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00478 sig68 sx[2] sx[6] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00477 vss u6.y0.xr2_x1_sig sig68 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00476 sig78 u1.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00475 vss rtl_map_7 sig81 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00474 sig77 sig81 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00473 sx[1] sig78 sig77 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00472 sig79 rtl_map_7 sx[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00471 vss u1.y0.xr2_x1_sig sig79 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00470 vss sig90 z[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00469 sig90 sx[10] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00468 vss vdd rtl_map_7 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00467 vss vdd rtl_map_9 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00466 sig95 u0.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00465 vss rtl_map_9 sig98 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00464 sig97 sig98 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00463 sx[0] sig95 sig97 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00462 sig94 rtl_map_9 sx[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00461 vss u0.y0.xr2_x1_sig sig94 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00460 vss sig110 cx[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00459 vss cx[2] sig146 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00458 sig146 u3.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00457 sig110 cx[2] sig147 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00456 sig147 u3.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00455 sig146 rtl_map_5 sig110 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00454 sig112 x[3] sig150 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00453 vss sig112 u3.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00452 sig150 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00451 vss sig119 cx[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00450 vss cx[1] sig157 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00449 sig157 u2.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00448 sig119 cx[1] sig158 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00447 sig158 u2.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00446 sig157 rtl_map_6 sig119 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00445 sig125 u2.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00444 vss cx[1] sig127 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00443 sig176 sig127 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00442 u2.y0.xr2_x1_sig sig125 sig176 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00441 sig171 cx[1] u2.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00440 vss u2.x1 sig171 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00439 vss vdd rtl_map_6 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00438 sig121 u2.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00437 vss rtl_map_6 sig123 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00436 sig166 sig123 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00435 sx[2] sig121 sig166 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00434 sig167 rtl_map_6 sx[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00433 vss u2.y0.xr2_x1_sig sig167 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00432 vss sig128 cx[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00431 vss cx[0] sig180 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00430 sig180 u1.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00429 sig128 cx[0] sig179 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00428 sig179 u1.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00427 sig180 rtl_map_7 sig128 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00426 sig137 x[0] sig193 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00425 vss sig137 u0.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00424 sig193 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00423 sig134 u1.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00422 vss cx[0] sig135 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00421 sig185 sig135 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00420 u1.y0.xr2_x1_sig sig134 sig185 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00419 sig186 cx[0] u1.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00418 vss u1.x1 sig186 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00417 sig143 u0.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00416 vss rtl_map_8 sig144 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00415 sig207 sig144 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00414 u0.y0.xr2_x1_sig sig143 sig207 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00413 sig201 rtl_map_8 u0.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00412 vss u0.x1 sig201 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00411 vss sig140 cx[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00410 vss rtl_map_8 sig198 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00409 sig198 u0.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00408 sig140 rtl_map_8 sig199 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00407 sig199 u0.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00406 sig198 rtl_map_9 sig140 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00405 sig155 u7.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00404 vss cx[6] sig156 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00403 sig151 sig156 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00402 u7.y0.xr2_x1_sig sig155 sig151 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00401 sig152 cx[6] u7.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00400 vss u7.x1 sig152 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00399 sig163 u7.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00398 vss sx[3] sig162 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00397 sig160 sig162 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00396 sx[7] sig163 sig160 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00395 sig161 sx[3] sx[7] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00394 vss u7.y0.xr2_x1_sig sig161 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00393 vss sig149 cx[7] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00392 vss cx[6] sig210 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00391 sig210 u7.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00390 sig149 cx[6] sig211 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00389 sig211 u7.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00388 sig210 sx[3] sig149 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00387 sig169 x[2] sig168 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00386 vss sig169 u2.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00385 sig168 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 sig175 x[1] sig173 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00383 vss sig175 u16.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 sig173 y[3] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 sig183 x[0] sig182 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 vss sig183 u15.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00379 sig182 y[3] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00378 sig165 x[1] sig164 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00377 vss sig165 u6.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00376 sig164 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00375 sig192 u15.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00374 vss rtl_map_1 sig190 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00373 sig187 sig190 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00372 u15.y0.xr2_x1_sig sig192 sig187 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00371 sig188 rtl_map_1 u15.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00370 vss u15.x1 sig188 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00369 vss sig184 cx[15] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00368 vss rtl_map_1 sig220 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00367 sig220 u15.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00366 sig184 rtl_map_1 sig218 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00365 sig218 u15.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00364 sig220 sx[11] sig184 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00363 vss vdd rtl_map_1 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00362 sig197 x[0] sig195 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00361 vss sig197 u20.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00360 sig195 y[4] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00359 sig205 u15.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00358 vss sx[11] sig206 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00357 sig202 sig206 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00356 sx[15] sig205 sig202 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00355 sig200 sx[11] sx[15] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00354 vss u15.y0.xr2_x1_sig sig200 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00353 sig178 x[1] sig177 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00352 vss sig178 u1.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00351 sig177 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00350 vss vdd rtl_map_8 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00349 vss sig209 z[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00348 sig209 sx[15] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00347 vss vdd rtl_map_0 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00346 sig232 x[2] sig271 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00345 vss sig232 u7.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00344 sig271 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00343 sig226 x[3] sig264 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00342 vss sig226 u8.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00341 sig264 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00340 sig228 u8.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00339 vss cx[7] sig231 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00338 sig266 sig231 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00337 u8.y0.xr2_x1_sig sig228 sig266 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00336 sig267 cx[7] u8.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00335 vss u8.x1 sig267 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 sig242 u16.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00333 vss cx[15] sig243 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00332 sig283 sig243 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00331 u16.y0.xr2_x1_sig sig242 sig283 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00330 sig284 cx[15] u16.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00329 vss u16.x1 sig284 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00328 vss sig237 cx[16] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00327 vss cx[15] sig277 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00326 sig277 u16.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00325 sig237 cx[15] sig278 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00324 sig278 u16.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00323 sig277 sx[12] sig237 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00322 sig233 x[1] sig272 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00321 vss sig233 u11.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00320 sig272 y[2] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00319 sig244 u16.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00318 vss sx[12] sig245 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00317 sig286 sig245 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00316 sx[16] sig244 sig286 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00315 sig285 sx[12] sx[16] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00314 vss u16.y0.xr2_x1_sig sig285 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00313 sig248 x[1] sig289 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00312 vss sig248 u21.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00311 sig289 y[4] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00310 vss sig252 cx[20] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00309 vss rtl_map_0 sig294 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00308 sig294 u20.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00307 sig252 rtl_map_0 sig291 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00306 sig291 u20.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00305 sig294 sx[16] sig252 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00304 sig255 u20.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00303 vss rtl_map_0 sig257 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00302 sig296 sig257 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 u20.y0.xr2_x1_sig sig255 sig296 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00300 sig295 rtl_map_0 u20.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00299 vss u20.x1 sig295 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00298 sig258 u20.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00297 vss sx[16] sig261 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00296 sig300 sig261 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 sx[20] sig258 sig300 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00294 sig299 sx[16] sx[20] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 vss u20.y0.xr2_x1_sig sig299 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 vss sig262 z[4] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 sig262 sx[20] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00290 vss sig306 cx[8] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 vss cx[7] sig307 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00288 sig307 u8.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00287 sig306 cx[7] sig308 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00286 sig308 u8.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00285 sig307 sx[4] sig306 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00284 sig268 u8.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00283 vss sx[4] sig269 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00282 sig314 sig269 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 sx[8] sig268 sig314 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 sig313 sx[4] sx[8] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00279 vss u8.y0.xr2_x1_sig sig313 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 sig276 u12.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00277 vss cx[11] sig273 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00276 sig317 sig273 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 u12.y0.xr2_x1_sig sig276 sig317 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 sig316 cx[11] u12.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00273 vss u12.x1 sig316 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00272 sig281 u12.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00271 vss sx[8] sig282 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00270 sig321 sig282 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00269 sx[12] sig281 sig321 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 sig319 sx[8] sx[12] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 vss u12.y0.xr2_x1_sig sig319 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00266 sig287 u11.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00265 vss cx[10] sig288 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00264 sig328 sig288 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00263 u11.y0.xr2_x1_sig sig287 sig328 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 sig327 cx[10] u11.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 vss u11.x1 sig327 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 vss sig322 cx[11] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00259 vss cx[10] sig324 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00258 sig324 u11.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00257 sig322 cx[10] sig323 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00256 sig323 u11.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00255 sig324 sx[7] sig322 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00254 sig292 u11.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00253 vss sx[7] sig293 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00252 sig332 sig293 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00251 sx[11] sig292 sig332 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00250 sig330 sx[7] sx[11] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00249 vss u11.y0.xr2_x1_sig sig330 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00248 sig297 u21.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00247 vss cx[20] sig298 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00246 sig341 sig298 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00245 u21.y0.xr2_x1_sig sig297 sig341 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 sig339 cx[20] u21.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 vss u21.x1 sig339 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00242 vss sig334 cx[21] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00241 vss cx[20] sig335 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00240 sig335 u21.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00239 sig334 cx[20] sig336 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00238 sig336 u21.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00237 sig335 sx[17] sig334 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00236 sig301 u21.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00235 vss sx[17] sig302 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00234 sig344 sig302 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00233 sx[21] sig301 sig344 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 sig342 sx[17] sx[21] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 vss u21.y0.xr2_x1_sig sig342 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 vss sig305 z[5] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 sig305 sx[21] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00228 vss vdd rtl_map_4 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00227 sig348 u4.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00226 vss rtl_map_4 sig351 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00225 sig385 sig351 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00224 sx[4] sig348 sig385 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00223 sig386 rtl_map_4 sx[4] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00222 vss u4.y0.xr2_x1_sig sig386 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00221 sig352 x[2] sig387 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 vss sig352 u12.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 sig387 y[2] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 vss sig356 cx[12] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 vss cx[11] sig389 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00216 sig389 u12.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00215 sig356 cx[11] sig388 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00214 sig388 u12.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00213 sig389 sx[8] sig356 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00212 sig357 x[2] sig390 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 vss sig357 u17.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00210 sig390 y[3] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00209 sig369 u17.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00208 vss sx[13] sig370 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00207 sig396 sig370 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 sx[17] sig369 sig396 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00205 sig395 sx[13] sx[17] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 vss u17.y0.xr2_x1_sig sig395 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00203 sig364 u17.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00202 vss cx[16] sig367 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00201 sig394 sig367 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 u17.y0.xr2_x1_sig sig364 sig394 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 sig393 cx[16] u17.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 vss u17.x1 sig393 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 vss sig361 cx[17] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 vss cx[16] sig392 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00195 sig392 u17.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00194 sig361 cx[16] sig391 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00193 sig391 u17.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00192 sig392 sx[13] sig361 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00191 sig371 x[2] sig397 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00190 vss sig371 u22.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00189 sig397 y[4] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00188 sig374 u22.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00187 vss cx[21] sig376 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00186 sig398 sig376 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00185 u22.y0.xr2_x1_sig sig374 sig398 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00184 sig399 cx[21] u22.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 vss u22.x1 sig399 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00182 vss sig383 z[6] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00181 sig383 sx[22] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00180 sig377 u22.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00179 vss sx[18] sig381 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00178 sig401 sig381 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00177 sx[22] sig377 sig401 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 sig400 sx[18] sx[22] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 vss u22.y0.xr2_x1_sig sig400 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 sig402 u4.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00173 vss cx[3] sig405 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00172 sig404 sig405 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 u4.y0.xr2_x1_sig sig402 sig404 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 sig403 cx[3] u4.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 vss u4.x1 sig403 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 vss sig408 cx[4] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 vss cx[3] sig409 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00166 sig409 u4.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00165 sig408 cx[3] sig407 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00164 sig407 u4.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00163 sig409 rtl_map_4 sig408 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00162 sig420 u13.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00161 vss sx[9] sig421 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00160 sig422 sig421 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 sx[13] sig420 sig422 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 sig419 sx[9] sx[13] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00157 vss u13.y0.xr2_x1_sig sig419 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00156 sig410 x[3] sig411 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00155 vss sig410 u13.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 sig411 y[2] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00153 sig414 u13.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00152 vss cx[12] sig415 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00151 sig418 sig415 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 u13.y0.xr2_x1_sig sig414 sig418 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 sig416 cx[12] u13.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00148 vss u13.x1 sig416 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 sig434 u18.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00146 vss cx[17] sig435 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00145 sig436 sig435 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00144 u18.y0.xr2_x1_sig sig434 sig436 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00143 sig432 cx[17] u18.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 vss u18.x1 sig432 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 sig430 x[3] sig431 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 vss sig430 u18.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 sig431 y[3] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 vss sig424 cx[18] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 vss cx[17] sig426 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00136 sig426 u18.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00135 sig424 cx[17] sig425 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00134 sig425 u18.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00133 sig426 sx[14] sig424 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00132 sig440 u18.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00131 vss sx[14] sig442 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00130 sig444 sig442 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 sx[18] sig440 sig444 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 sig443 sx[14] sx[18] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00127 vss u18.y0.xr2_x1_sig sig443 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 vss sig437 cx[22] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 vss cx[21] sig438 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00124 sig438 u22.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00123 sig437 cx[21] sig439 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00122 sig439 u22.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00121 sig438 sx[18] sig437 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00120 vss sig446 z[7] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 sig446 sx[23] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00118 sig455 x[4] sig507 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 vss sig455 u4.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 sig507 y[0] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 sig451 u9.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00114 vss cx[8] sig454 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00113 sig505 sig454 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 u9.y0.xr2_x1_sig sig451 sig505 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 sig506 cx[8] u9.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 vss u9.x1 sig506 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 sig459 u9.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00108 vss cx[4] sig461 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 sig508 sig461 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 sx[9] sig459 sig508 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 sig509 cx[4] sx[9] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 vss u9.y0.xr2_x1_sig sig509 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 sig466 x[4] sig512 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 vss sig466 u19.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 sig512 y[3] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 vss sig463 cx[13] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 vss cx[12] sig511 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00098 sig511 u13.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00097 sig463 cx[12] sig510 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00096 sig510 u13.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00095 sig511 sx[9] sig463 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00094 vss sig472 cx[19] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 vss cx[18] sig514 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00092 sig514 u19.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00091 sig472 cx[18] sig513 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00090 sig513 u19.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00089 sig514 cx[14] sig472 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00088 sig480 u19.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00087 vss cx[14] sig483 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00086 sig518 sig483 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 sx[19] sig480 sig518 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00084 sig517 cx[14] sx[19] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 vss u19.y0.xr2_x1_sig sig517 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 sig478 u19.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00081 vss cx[18] sig479 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00080 sig515 sig479 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 u19.y0.xr2_x1_sig sig478 sig515 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 sig516 cx[18] u19.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 vss u19.x1 sig516 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 sig487 x[4] sig519 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00075 vss sig487 u24.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 sig519 y[4] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 sig488 x[3] sig520 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 vss sig488 u23.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 sig520 y[4] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 sig497 u23.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 vss cx[22] sig499 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00068 sig524 sig499 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 u23.y0.xr2_x1_sig sig497 sig524 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 sig523 cx[22] u23.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 vss u23.x1 sig523 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 vss sig495 cx[23] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 vss cx[22] sig522 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00062 sig522 u23.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00061 sig495 cx[22] sig521 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00060 sig521 u23.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00059 sig522 sx[19] sig495 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00058 sig501 u23.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00057 vss sx[19] sig503 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 sig526 sig503 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 sx[23] sig501 sig526 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 sig525 sx[19] sx[23] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 vss u23.y0.xr2_x1_sig sig525 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 vss sig530 cx[9] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 vss cx[8] sig531 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00050 sig531 u9.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00049 sig530 cx[8] sig532 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00048 sig532 u9.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00047 sig531 cx[4] sig530 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00046 sig528 x[4] sig529 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 vss sig528 u9.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 sig529 y[1] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 sig536 x[4] sig534 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 vss sig536 u14.x1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 sig534 y[2] vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 sig540 u14.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00039 vss cx[13] sig544 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 sig543 sig544 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 u14.y0.xr2_x1_sig sig540 sig543 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 sig541 cx[13] u14.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 vss u14.x1 sig541 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 sig546 u14.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 vss cx[9] sig548 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 sig545 sig548 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 sx[14] sig546 sig545 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 sig547 cx[9] sx[14] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 vss u14.y0.xr2_x1_sig sig547 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 vss sig537 cx[14] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 vss cx[13] sig538 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00026 sig538 u14.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00025 sig537 cx[13] sig539 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00024 sig539 u14.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00023 sig538 cx[9] sig537 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00022 vss sig560 cx[24] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 vss cx[23] sig559 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00020 sig559 u24.x1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00019 sig560 cx[23] sig561 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00018 sig561 u24.x1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00017 sig559 cx[19] sig560 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00016 sig556 u24.x1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 vss cx[23] sig557 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 sig558 sig557 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 u24.y0.xr2_x1_sig sig556 sig558 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 sig555 cx[23] u24.y0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 vss u24.x1 sig555 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 vss sig563 z[8] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 sig563 sx[24] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00008 vss sig565 z[9] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 sig565 cx[24] vss vss tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00006 sig549 u24.y0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 vss cx[19] sig552 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 sig551 sig552 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 sx[24] sig549 sig551 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 sig553 cx[19] sx[24] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 vss u24.y0.xr2_x1_sig sig553 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C576 sig576 vss 8.58e-15
C574 sig574 vss 9.7e-15
C573 sig573 vss 9.7e-15
C572 sig572 vss 9.7e-15
C571 sig571 vss 9.7e-15
C569 sig569 vss 8.58e-15
C568 sig568 vss 8.58e-15
C565 sig565 vss 1.568e-14
C564 z[9] vss 2.659e-14
C563 sig563 vss 1.568e-14
C562 cx[24] vss 6.053e-14
C560 sig560 vss 2.299e-14
C559 sig559 vss 4.11e-15
C557 sig557 vss 2.596e-14
C556 sig556 vss 2.16e-14
C554 sx[24] vss 8.739e-14
C552 sig552 vss 2.596e-14
C550 u24.y0.xr2_x1_sig vss 6.351e-14
C549 sig549 vss 2.16e-14
C548 sig548 vss 2.596e-14
C546 sig546 vss 2.16e-14
C544 sig544 vss 2.596e-14
C542 u14.y0.xr2_x1_sig vss 5.991e-14
C540 sig540 vss 2.16e-14
C538 sig538 vss 4.11e-15
C537 sig537 vss 2.299e-14
C536 sig536 vss 1.8635e-14
C535 u14.x1 vss 1.0771e-13
C533 cx[9] vss 1.1845e-13
C531 sig531 vss 4.11e-15
C530 sig530 vss 2.299e-14
C528 sig528 vss 1.8635e-14
C527 z[8] vss 4.387e-14
C522 sig522 vss 4.11e-15
C514 sig514 vss 4.11e-15
C511 sig511 vss 4.11e-15
C503 sig503 vss 2.596e-14
C502 sig502 vss 9.7e-15
C501 sig501 vss 2.16e-14
C500 sig500 vss 9.7e-15
C499 sig499 vss 2.596e-14
C498 u23.y0.xr2_x1_sig vss 5.751e-14
C497 sig497 vss 2.16e-14
C496 sig496 vss 9.7e-15
C495 sig495 vss 2.299e-14
C494 cx[23] vss 1.0376e-13
C491 sig491 vss 8.58e-15
C490 sig490 vss 8.58e-15
C489 u23.x1 vss 1.0291e-13
C488 sig488 vss 1.8635e-14
C487 sig487 vss 1.8635e-14
C486 u24.x1 vss 1.1915e-13
C485 sig485 vss 9.7e-15
C484 sx[19] vss 1.2419e-13
C483 sig483 vss 2.596e-14
C482 sig482 vss 9.7e-15
C480 sig480 vss 2.16e-14
C479 sig479 vss 2.596e-14
C478 sig478 vss 2.16e-14
C477 u19.y0.xr2_x1_sig vss 5.751e-14
C476 sig476 vss 9.7e-15
C475 sig475 vss 8.58e-15
C474 cx[14] vss 1.1653e-13
C472 sig472 vss 2.299e-14
C471 cx[19] vss 1.2373e-13
C470 sig470 vss 8.58e-15
C469 u19.x1 vss 1.0291e-13
C468 sig468 vss 9.7e-15
C467 cx[13] vss 1.1456e-13
C466 sig466 vss 1.8635e-14
C465 sig465 vss 9.7e-15
C464 sig464 vss 8.58e-15
C463 sig463 vss 2.299e-14
C461 sig461 vss 2.596e-14
C460 sig460 vss 9.7e-15
C459 sig459 vss 2.16e-14
C457 x[4] vss 1.9162e-13
C456 sig456 vss 8.58e-15
C455 sig455 vss 1.8635e-14
C454 sig454 vss 2.596e-14
C453 u9.x1 vss 1.0819e-13
C452 u9.y0.xr2_x1_sig vss 6.711e-14
C451 sig451 vss 2.16e-14
C450 sig450 vss 9.7e-15
C449 sig449 vss 9.7e-15
C447 sx[23] vss 5.979e-14
C446 sig446 vss 1.568e-14
C445 z[7] vss 2.371e-14
C442 sig442 vss 2.596e-14
C441 cx[22] vss 1.2104e-13
C440 sig440 vss 2.16e-14
C438 sig438 vss 4.11e-15
C437 sig437 vss 2.299e-14
C435 sig435 vss 2.596e-14
C434 sig434 vss 2.16e-14
C433 u18.y0.xr2_x1_sig vss 7.311e-14
C430 sig430 vss 1.8635e-14
C429 cx[18] vss 1.1944e-13
C428 u18.x1 vss 1.1131e-13
C427 sx[14] vss 1.4459e-13
C426 sig426 vss 4.11e-15
C424 sig424 vss 2.299e-14
C423 sx[9] vss 1.1987e-13
C421 sig421 vss 2.596e-14
C420 sig420 vss 2.16e-14
C417 u13.y0.xr2_x1_sig vss 5.991e-14
C415 sig415 vss 2.596e-14
C414 sig414 vss 2.16e-14
C413 u13.x1 vss 1.0627e-13
C412 cx[4] vss 1.1389e-13
C410 sig410 vss 1.8635e-14
C409 sig409 vss 4.11e-15
C408 sig408 vss 2.299e-14
C406 u4.x1 vss 1.1803e-13
C405 sig405 vss 2.596e-14
C402 sig402 vss 2.16e-14
C392 sig392 vss 4.11e-15
C389 sig389 vss 4.11e-15
C383 sig383 vss 1.568e-14
C382 z[6] vss 2.371e-14
C381 sig381 vss 2.596e-14
C380 sx[18] vss 1.0587e-13
C379 sx[22] vss 5.619e-14
C378 sig378 vss 9.7e-15
C377 sig377 vss 2.16e-14
C376 sig376 vss 2.596e-14
C375 u22.y0.xr2_x1_sig vss 5.991e-14
C374 sig374 vss 2.16e-14
C373 sig373 vss 9.7e-15
C372 u22.x1 vss 1.1227e-13
C371 sig371 vss 1.8635e-14
C370 sig370 vss 2.596e-14
C369 sig369 vss 2.16e-14
C368 sig368 vss 9.7e-15
C367 sig367 vss 2.596e-14
C366 u17.y0.xr2_x1_sig vss 5.991e-14
C365 cx[17] vss 1.2824e-13
C364 sig364 vss 2.16e-14
C363 sig363 vss 9.7e-15
C362 sx[13] vss 1.1291e-13
C361 sig361 vss 2.299e-14
C359 sig359 vss 8.58e-15
C358 u17.x1 vss 1.0771e-13
C357 sig357 vss 1.8635e-14
C356 sig356 vss 2.299e-14
C355 cx[12] vss 1.256e-13
C353 sig353 vss 8.58e-15
C352 sig352 vss 1.8635e-14
C351 sig351 vss 2.596e-14
C350 u4.y0.xr2_x1_sig vss 5.751e-14
C349 rtl_map_4 vss 9.269e-14
C348 sig348 vss 2.16e-14
C347 sig347 vss 9.7e-15
C346 z[5] vss 2.371e-14
C345 sig345 vss 9.7e-15
C343 sx[21] vss 5.619e-14
C340 sig340 vss 9.7e-15
C338 cx[21] vss 1.232e-13
C335 sig335 vss 4.11e-15
C334 sig334 vss 2.299e-14
C333 sig333 vss 8.58e-15
C331 sig331 vss 9.7e-15
C329 sig329 vss 9.7e-15
C325 sig325 vss 8.58e-15
C324 sig324 vss 4.11e-15
C322 sig322 vss 2.299e-14
C320 sig320 vss 9.7e-15
C318 sig318 vss 9.7e-15
C315 sig315 vss 9.7e-15
C312 cx[8] vss 1.468e-13
C310 sig310 vss 8.58e-15
C307 sig307 vss 4.11e-15
C306 sig306 vss 2.299e-14
C305 sig305 vss 1.568e-14
C304 sx[17] vss 1.2059e-13
C303 u21.y0.xr2_x1_sig vss 5.751e-14
C302 sig302 vss 2.596e-14
C301 sig301 vss 2.16e-14
C298 sig298 vss 2.596e-14
C297 sig297 vss 2.16e-14
C294 sig294 vss 4.11e-15
C293 sig293 vss 2.596e-14
C292 sig292 vss 2.16e-14
C290 u11.y0.xr2_x1_sig vss 5.991e-14
C288 sig288 vss 2.596e-14
C287 sig287 vss 2.16e-14
C282 sig282 vss 2.596e-14
C281 sig281 vss 2.16e-14
C280 sx[8] vss 1.1867e-13
C279 u12.y0.xr2_x1_sig vss 5.991e-14
C277 sig277 vss 4.11e-15
C276 sig276 vss 2.16e-14
C275 cx[11] vss 1.3552e-13
C274 u12.x1 vss 1.0675e-13
C273 sig273 vss 2.596e-14
C270 sx[4] vss 1.0211e-13
C269 sig269 vss 2.596e-14
C268 sig268 vss 2.16e-14
C263 z[4] vss 2.371e-14
C262 sig262 vss 1.568e-14
C261 sig261 vss 2.596e-14
C260 sig260 vss 9.7e-15
C259 sx[20] vss 5.619e-14
C258 sig258 vss 2.16e-14
C257 sig257 vss 2.596e-14
C256 u20.y0.xr2_x1_sig vss 5.751e-14
C255 sig255 vss 2.16e-14
C254 sig254 vss 9.7e-15
C252 sig252 vss 2.299e-14
C251 cx[20] vss 1.1264e-13
C250 u21.x1 vss 1.1443e-13
C249 sig249 vss 8.58e-15
C248 sig248 vss 1.8635e-14
C247 sx[16] vss 1.2131e-13
C246 sig246 vss 9.7e-15
C245 sig245 vss 2.596e-14
C244 sig244 vss 2.16e-14
C243 sig243 vss 2.596e-14
C242 sig242 vss 2.16e-14
C241 sig241 vss 9.7e-15
C240 u16.y0.xr2_x1_sig vss 5.991e-14
C239 cx[16] vss 1.3304e-13
C238 sx[12] vss 1.1291e-13
C237 sig237 vss 2.299e-14
C235 sig235 vss 8.58e-15
C234 u11.x1 vss 1.2859e-13
C233 sig233 vss 1.8635e-14
C232 sig232 vss 1.8635e-14
C231 sig231 vss 2.596e-14
C230 sig230 vss 9.7e-15
C229 u8.y0.xr2_x1_sig vss 5.991e-14
C228 sig228 vss 2.16e-14
C227 u8.x1 vss 1.1123e-13
C226 sig226 vss 1.8635e-14
C225 sig225 vss 9.7e-15
C224 rtl_map_0 vss 1.1496e-13
C223 sig223 vss 9.7e-15
C222 cx[15] vss 1.4024e-13
C220 sig220 vss 4.11e-15
C219 sig219 vss 8.58e-15
C217 sig217 vss 9.7e-15
C216 sig216 vss 9.7e-15
C215 cx[7] vss 1.2704e-13
C212 sig212 vss 8.58e-15
C210 sig210 vss 4.11e-15
C209 sig209 vss 1.568e-14
C208 z[3] vss 2.371e-14
C206 sig206 vss 2.596e-14
C205 sig205 vss 2.16e-14
C204 sx[11] vss 1.3331e-13
C203 sx[15] vss 5.979e-14
C198 sig198 vss 4.11e-15
C197 sig197 vss 1.8635e-14
C196 y[4] vss 2.7149e-13
C194 u20.x1 vss 1.0771e-13
C192 sig192 vss 2.16e-14
C191 rtl_map_1 vss 1.0392e-13
C190 sig190 vss 2.596e-14
C189 u15.y0.xr2_x1_sig vss 6.711e-14
C184 sig184 vss 2.299e-14
C183 sig183 vss 1.8635e-14
C181 u15.x1 vss 1.0651e-13
C180 sig180 vss 4.11e-15
C178 sig178 vss 1.8635e-14
C175 sig175 vss 1.8635e-14
C174 y[3] vss 3.0277e-13
C172 u16.x1 vss 1.1443e-13
C170 x[2] vss 2.4538e-13
C169 sig169 vss 1.8635e-14
C165 sig165 vss 1.8635e-14
C163 sig163 vss 2.16e-14
C162 sig162 vss 2.596e-14
C159 sx[7] vss 1.4819e-13
C157 sig157 vss 4.11e-15
C156 sig156 vss 2.596e-14
C155 sig155 vss 2.16e-14
C154 u7.x1 vss 1.2091e-13
C153 u7.y0.xr2_x1_sig vss 5.991e-14
C149 sig149 vss 2.299e-14
C148 x[1] vss 2.0586e-13
C146 sig146 vss 4.11e-15
C144 sig144 vss 2.596e-14
C143 sig143 vss 2.16e-14
C142 sig142 vss 9.7e-15
C141 rtl_map_8 vss 1.1304e-13
C140 sig140 vss 2.299e-14
C138 sig138 vss 8.58e-15
C137 sig137 vss 1.8635e-14
C136 u0.x1 vss 1.0531e-13
C135 sig135 vss 2.596e-14
C134 sig134 vss 2.16e-14
C133 sig133 vss 9.7e-15
C131 u1.x1 vss 1.1491e-13
C130 cx[0] vss 1.3528e-13
C129 sig129 vss 8.58e-15
C128 sig128 vss 2.299e-14
C127 sig127 vss 2.596e-14
C126 sig126 vss 9.7e-15
C125 sig125 vss 2.16e-14
C124 sig124 vss 9.7e-15
C123 sig123 vss 2.596e-14
C122 u2.y0.xr2_x1_sig vss 6.351e-14
C121 sig121 vss 2.16e-14
C120 cx[1] vss 1.3904e-13
C119 sig119 vss 2.299e-14
C117 u2.x1 vss 1.2083e-13
C116 rtl_map_6 vss 9.341e-14
C115 sig115 vss 8.58e-15
C114 y[0] vss 3.4405e-13
C113 x[3] vss 2.6938e-13
C112 sig112 vss 1.8635e-14
C111 cx[3] vss 1.5176e-13
C110 sig110 vss 2.299e-14
C108 sig108 vss 8.58e-15
C107 sig107 vss 9.7e-15
C106 sig106 vss 9.7e-15
C105 sig105 vss 9.7e-15
C104 sig104 vss 9.7e-15
C103 sig103 vss 9.7e-15
C101 sig101 vss 8.58e-15
C100 sig100 vss 9.7e-15
C99 sig99 vss 9.7e-15
C98 sig98 vss 2.596e-14
C96 u0.y0.xr2_x1_sig vss 6.231e-14
C95 sig95 vss 2.16e-14
C93 rtl_map_9 vss 9.517e-14
C91 z[2] vss 5.707e-14
C90 sig90 vss 1.568e-14
C88 sx[10] vss 5.859e-14
C86 sig86 vss 2.596e-14
C84 sig84 vss 2.16e-14
C81 sig81 vss 2.596e-14
C80 u1.y0.xr2_x1_sig vss 6.951e-14
C78 sig78 vss 2.16e-14
C76 rtl_map_7 vss 8.909e-14
C73 sig73 vss 4.11e-15
C71 sig71 vss 2.596e-14
C69 sig69 vss 2.16e-14
C66 u6.y0.xr2_x1_sig vss 5.991e-14
C64 sig64 vss 2.596e-14
C63 sig63 vss 4.11e-15
C62 cx[6] vss 1.4264e-13
C61 sig61 vss 2.16e-14
C59 sx[2] vss 1.2371e-13
C57 sig57 vss 2.299e-14
C56 sig56 vss 4.11e-15
C53 u6.x1 vss 1.1971e-13
C52 cx[2] vss 1.34e-13
C50 sig50 vss 2.596e-14
C48 u3.x1 vss 1.1419e-13
C47 sig47 vss 2.16e-14
C45 sig45 vss 2.596e-14
C44 u3.y0.xr2_x1_sig vss 6.351e-14
C42 sx[3] vss 1.2491e-13
C40 sig40 vss 2.16e-14
C39 vss vss 6.36869e-12
C38 sx[0] vss 5.859e-14
C37 sig37 vss 1.568e-14
C36 z[0] vss 2.659e-14
C35 sig35 vss 1.568e-14
C34 z[1] vss 4.387e-14
C33 sig33 vss 2.596e-14
C32 sig32 vss 2.16e-14
C31 sx[5] vss 5.859e-14
C30 sig30 vss 9.7e-15
C29 sig29 vss 2.596e-14
C28 u10.y0.xr2_x1_sig vss 6.111e-14
C27 sig27 vss 9.7e-15
C26 sig26 vss 2.16e-14
C25 cx[10] vss 1.7144e-13
C24 rtl_map_2 vss 1.1744e-13
C23 sx[6] vss 1.2659e-13
C22 sig22 vss 2.299e-14
C20 y[2] vss 3.4597e-13
C19 sig19 vss 8.58e-15
C18 u10.x1 vss 1.0771e-13
C17 sig17 vss 1.8635e-14
C16 sx[1] vss 1.5803e-13
C15 sig15 vss 2.299e-14
C14 cx[5] vss 1.1504e-13
C12 sig12 vss 8.58e-15
C11 u5.y0.xr2_x1_sig vss 1.2111e-13
C10 sig10 vss 9.7e-15
C9 sig9 vss 2.596e-14
C8 sig8 vss 2.16e-14
C7 rtl_map_3 vss 1.2232e-13
C6 x[0] vss 2.5402e-13
C5 y[1] vss 3.4717e-13
C4 u5.x1 vss 1.2907e-13
C3 sig3 vss 1.8635e-14
C2 rtl_map_5 vss 9.749e-14
C1 vdd vss 6.61006e-12
.ends mul5b_cougar

