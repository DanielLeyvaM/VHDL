* Spice description of mul2b_cougar
* Spice driver version -1208873308
* Date ( dd/mm/yyyy hh:mm:ss ): 28/10/2020 at 14:06:10

* INTERF vdd vss x[0] x[1] y[0] y[1] z[0] z[1] z[2] z[3] 


.subckt mul2b_cougar 31 18 27 26 28 23 21 7 24 3 
* NET 3 = z[3]
* NET 7 = z[1]
* NET 12 = aux2
* NET 17 = aux1
* NET 18 = vss
* NET 21 = z[0]
* NET 22 = inv_x2_sig
* NET 23 = y[1]
* NET 24 = z[2]
* NET 26 = x[1]
* NET 27 = x[0]
* NET 28 = y[0]
* NET 29 = not_aux0
* NET 31 = vdd
Mtr_00050 31 22 25 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 24 25 31 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00048 31 23 25 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 25 26 31 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 29 30 31 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00045 31 28 30 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 30 27 31 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 22 29 31 31 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00042 21 20 31 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00041 31 29 20 31 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00040 17 16 31 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00039 31 28 16 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 16 26 31 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 12 11 31 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00036 31 23 11 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 11 27 31 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 8 12 31 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 31 17 9 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 7 8 1 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00031 1 17 31 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00030 1 9 7 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00029 31 12 1 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00028 3 2 31 31 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00027 31 17 2 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 2 12 31 31 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 18 25 24 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 13 22 18 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 14 26 13 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 25 23 14 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 30 27 19 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 18 30 29 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 19 28 18 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 18 29 22 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 18 20 21 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 20 29 18 18 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00015 16 26 15 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 18 16 17 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 15 28 18 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 11 27 10 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 18 11 12 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 10 23 18 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 9 17 18 18 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 18 12 8 18 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 6 8 18 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 7 9 6 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 5 12 7 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 18 17 5 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 2 12 4 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 18 2 3 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 4 17 18 18 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C32 1 18 9.7e-15
C30 2 18 1.8635e-14
C29 3 18 2.371e-14
C25 7 18 4.537e-14
C24 8 18 2.596e-14
C23 9 18 2.16e-14
C21 11 18 1.8635e-14
C20 12 18 8.2e-14
C16 16 18 1.8635e-14
C15 17 18 1.0506e-13
C14 18 18 3.2572e-13
C12 20 18 1.568e-14
C11 21 18 2.539e-14
C10 22 18 4.959e-14
C9 23 18 7.455e-14
C8 24 18 5.235e-14
C7 25 18 2.605e-14
C6 26 18 5.915e-14
C5 27 18 6.009e-14
C4 28 18 6.789e-14
C3 29 18 9.168e-14
C2 30 18 1.8635e-14
C1 31 18 3.4392e-13
.ends mul2b_cougar

