* Spice description of act5_cougar
* Spice driver version -1208955228
* Date ( dd/mm/yyyy hh:mm:ss ): 22/11/2020 at 11:54:04

* INTERF clk ctrl ctrl1 dh[0] dh[1] dh[2] dh[3] dm[0] dm[1] dm[2] dm[3] rst 
* INTERF uh[0] uh[1] uh[2] uh[3] um[0] um[1] um[2] um[3] vdd vss 


.subckt act5_cougar 1810 1244 184 839 476 186 22 1228 1157 1061 949 1708 846 845 841 479 1728 1607 1474 1345 1814 1727 
* NET 22 = dh[3]
* NET 24 = cdm_0_ins.sff_s
* NET 28 = cdm_0_ins.y
* NET 30 = cdm_0_ins.sff_m
* NET 32 = cdm_0_ins.u
* NET 33 = cdm_0_ins.nckr
* NET 34 = cdm_0_ins.ckr
* NET 39 = xr2_x1_2_sig
* NET 41 = on12_x1_4_sig
* NET 42 = noa22_x1_13_sig
* NET 45 = a3_x2_2_sig
* NET 48 = na2_x1_10_sig
* NET 54 = stop
* NET 56 = stop_ins.sff_s
* NET 57 = stop_ins.y
* NET 59 = stop_ins.sff_m
* NET 61 = stop_ins.u
* NET 62 = stop_ins.ckr
* NET 63 = stop_ins.nckr
* NET 65 = inv_x2_4_sig
* NET 70 = noa22_x1_6_sig
* NET 73 = on12_x1_sig
* NET 75 = cdh_2_ins.y
* NET 77 = cdh_2_ins.sff_m
* NET 78 = cdh_2_ins.sff_s
* NET 79 = noa22_x1_5_sig
* NET 81 = cdh_2_ins.nckr
* NET 82 = cdh_2_ins.u
* NET 83 = cdh_2_ins.ckr
* NET 85 = cdm_1_ins.y
* NET 86 = cdm_1_ins.sff_s
* NET 87 = cdm_1_ins.u
* NET 88 = cdm_1_ins.sff_m
* NET 91 = cdm_1_ins.ckr
* NET 92 = cdm_1_ins.nckr
* NET 95 = a2_x2_5_sig
* NET 96 = ao22_x2_sig
* NET 101 = a3_x2_3_sig
* NET 102 = an12_x1_2_sig
* NET 105 = aux60
* NET 108 = oa22_x2_11_sig
* NET 112 = na2_x1_11_sig
* NET 114 = cdh_0_ins.sff_s
* NET 115 = cdh_0_ins.y
* NET 118 = cdh_0_ins.sff_m
* NET 119 = cdh_0_ins.u
* NET 120 = cdh_0_ins.ckr
* NET 121 = cdh_0_ins.nckr
* NET 122 = inv_x2_3_sig
* NET 125 = noa22_x1_3_sig
* NET 127 = noa22_x1_2_sig
* NET 128 = oa22_x2_sig
* NET 132 = inv_x2_2_sig
* NET 134 = noa22_x1_sig
* NET 138 = a2_x2_7_sig
* NET 141 = oa22_x2_15_sig
* NET 145 = cum_0_ins.sff_s
* NET 146 = noa22_x1_16_sig
* NET 147 = cum_0_ins.y
* NET 149 = cum_0_ins.u
* NET 150 = cum_0_ins.sff_m
* NET 152 = cum_0_ins.nckr
* NET 153 = cum_0_ins.ckr
* NET 155 = mbk_buf_not_aux128
* NET 158 = xr2_x1_sig
* NET 166 = nxr2_x1_sig
* NET 184 = ctrl1
* NET 186 = dh[2]
* NET 190 = cdm_3_ins.y
* NET 192 = cdm_3_ins.sff_m
* NET 193 = cdm_3_ins.sff_s
* NET 194 = cdm_3_ins.u
* NET 196 = cdm_3_ins.ckr
* NET 197 = cdm_3_ins.nckr
* NET 198 = noa22_x1_15_sig
* NET 202 = oa2ao222_x2_sig
* NET 203 = inv_x2_7_sig
* NET 212 = no4_x1_5_sig
* NET 213 = a2_x2_6_sig
* NET 215 = aux63
* NET 216 = oa22_x2_2_sig
* NET 219 = na2_x1_6_sig
* NET 223 = no4_x1_2_sig
* NET 224 = aux32
* NET 226 = nao22_x1_sig
* NET 229 = aux4
* NET 230 = not_aux4
* NET 233 = oa22_x2_4_sig
* NET 236 = not_aux128
* NET 238 = a2_x2_2_sig
* NET 244 = maquina_ins.y
* NET 246 = maquina_ins.sff_m
* NET 247 = maquina_ins.sff_s
* NET 248 = no2_x1_sig
* NET 250 = maquina_ins.nckr
* NET 251 = maquina_ins.u
* NET 252 = maquina_ins.ckr
* NET 256 = rtlalc_9_2_ins.u
* NET 258 = rtlalc_9_2_ins.ckr
* NET 259 = rtlalc_9_2_ins.nckr
* NET 265 = not_aux44
* NET 267 = aux61
* NET 268 = aux62
* NET 272 = not_aux62
* NET 279 = na2_x1_3_sig
* NET 282 = na2_x1_4_sig
* NET 296 = cdh_1_ins.u
* NET 297 = cdh_1_ins.ckr
* NET 298 = cdh_1_ins.nckr
* NET 300 = rtlalc_9[2]
* NET 301 = rtlalc_9_2_ins.sff_s
* NET 302 = rtlalc_9_2_ins.sff_m
* NET 303 = rtlalc_9_2_ins.y
* NET 309 = oa22_x2_14_sig
* NET 312 = na3_x1_11_sig
* NET 315 = o3_x2_9_sig
* NET 319 = not_aux67
* NET 326 = o3_x2_8_sig
* NET 333 = not_aux24
* NET 337 = mbk_buf_aux4
* NET 341 = na4_x1_3_sig
* NET 344 = o4_x2_3_sig
* NET 346 = mbk_buf_not_aux3
* NET 347 = na3_x1_3_sig
* NET 350 = not_cdh[3]
* NET 351 = not_aux18
* NET 361 = na3_x1_5_sig
* NET 363 = noa22_x1_4_sig
* NET 365 = cdh_1_ins.sff_s
* NET 367 = cdh_1_ins.sff_m
* NET 368 = cdh_1_ins.y
* NET 373 = cdm_2_ins.y
* NET 374 = cdm_2_ins.sff_s
* NET 376 = cdm_2_ins.u
* NET 377 = cdm_2_ins.sff_m
* NET 380 = na2_x1_13_sig
* NET 381 = cdm_2_ins.nckr
* NET 382 = cdm_2_ins.ckr
* NET 384 = an12_x1_3_sig
* NET 386 = aux64
* NET 391 = oa22_x2_12_sig
* NET 392 = o4_x2_sig
* NET 395 = oa22_x2_13_sig
* NET 396 = noa22_x1_14_sig
* NET 398 = na2_x1_12_sig
* NET 399 = a3_x2_4_sig
* NET 400 = not_aux59
* NET 402 = o2_x2_5_sig
* NET 406 = cuh_2_ins.sff_s
* NET 407 = cuh_2_ins.y
* NET 409 = cuh_2_ins.sff_m
* NET 411 = cuh_2_ins.u
* NET 412 = cuh_2_ins.ckr
* NET 413 = cuh_2_ins.nckr
* NET 414 = na3_x1_4_sig
* NET 415 = not_aux118
* NET 417 = na3_x1_2_sig
* NET 420 = na2_x1_2_sig
* NET 421 = o2_x2_2_sig
* NET 424 = not_aux3
* NET 430 = cdh_3_ins.sff_s
* NET 431 = cdh_3_ins.y
* NET 433 = cdh_3_ins.sff_m
* NET 434 = cdh_3_ins.nckr
* NET 435 = cdh_3_ins.u
* NET 436 = cdh_3_ins.ckr
* NET 438 = noa22_x1_7_sig
* NET 439 = na3_x1_7_sig
* NET 440 = oa22_x2_5_sig
* NET 441 = o3_x2_2_sig
* NET 444 = na3_x1_6_sig
* NET 445 = not_aux25
* NET 446 = oa22_x2_3_sig
* NET 476 = dh[1]
* NET 479 = uh[3]
* NET 482 = on12_x1_5_sig
* NET 484 = o4_x2_2_sig
* NET 488 = not_cdm[0]
* NET 489 = not_aux45
* NET 498 = o2_x2_3_sig
* NET 501 = oa22_x2_8_sig
* NET 502 = na3_x1_10_sig
* NET 503 = noa22_x1_10_sig
* NET 506 = not_aux54
* NET 508 = a4_x2_sig
* NET 514 = not_aux16
* NET 519 = na2_x1_5_sig
* NET 521 = mbk_buf_not_aux4
* NET 522 = an12_x1_sig
* NET 523 = no4_x1_sig
* NET 526 = a4_x2_2_sig
* NET 532 = rtlalc_9[1]
* NET 533 = rtlalc_9_1_ins.y
* NET 534 = rtlalc_9_1_ins.sff_s
* NET 536 = rtlalc_9_1_ins.u
* NET 538 = rtlalc_9_1_ins.sff_m
* NET 541 = rtlalc_9_1_ins.ckr
* NET 542 = rtlalc_9_1_ins.nckr
* NET 549 = mbk_buf_not_aux1
* NET 551 = o2_x2_sig
* NET 553 = not_cdh[1]
* NET 554 = o3_x2_3_sig
* NET 557 = inv_x2_5_sig
* NET 559 = aux114
* NET 560 = not_aux31
* NET 561 = o3_x2_sig
* NET 564 = rtlalc_9[3]
* NET 566 = rtlalc_9_3_ins.sff_s
* NET 567 = rtlalc_9_3_ins.y
* NET 569 = rtlalc_9_3_ins.u
* NET 571 = rtlalc_9_3_ins.sff_m
* NET 572 = rtlalc_9_3_ins.nckr
* NET 573 = rtlalc_9_3_ins.ckr
* NET 574 = no2_x1_3_sig
* NET 576 = not_aux33
* NET 578 = na4_x1_2_sig
* NET 580 = aux33
* NET 582 = o3_x2_6_sig
* NET 587 = ao2o22_x2_3_sig
* NET 588 = cdh[2]
* NET 595 = not_cuh[2]
* NET 596 = not_cdm[2]
* NET 598 = no4_x1_4_sig
* NET 601 = not_aux37
* NET 602 = not_cdh[0]
* NET 606 = ao2o22_x2_4_sig
* NET 610 = not_aux41
* NET 611 = not_cdh[2]
* NET 612 = cdh[3]
* NET 617 = ao2o22_x2_2_sig
* NET 618 = cdh[1]
* NET 622 = not_aux14
* NET 623 = na2_x1_14_sig
* NET 625 = na2_x1_15_sig
* NET 626 = a3_x2_6_sig
* NET 628 = no2_x1_4_sig
* NET 631 = cum_3_ins.sff_s
* NET 632 = cum_3_ins.y
* NET 634 = cum_3_ins.sff_m
* NET 635 = noa22_x1_17_sig
* NET 637 = cum_3_ins.u
* NET 638 = cum_3_ins.ckr
* NET 639 = cum_3_ins.nckr
* NET 660 = cuh_1_ins.sff_s
* NET 662 = cuh_1_ins.y
* NET 664 = cuh_1_ins.u
* NET 666 = cuh_1_ins.sff_m
* NET 670 = not_aux32
* NET 671 = cuh_1_ins.ckr
* NET 672 = cuh_1_ins.nckr
* NET 673 = noa22_x1_9_sig
* NET 675 = na3_x1_9_sig
* NET 679 = oa22_x2_7_sig
* NET 681 = not_aux115
* NET 682 = not_aux48
* NET 683 = o3_x2_5_sig
* NET 685 = not_cdm[1]
* NET 690 = on12_x1_3_sig
* NET 693 = no2_x1_2_sig
* NET 694 = na2_x1_9_sig
* NET 695 = o3_x2_7_sig
* NET 701 = o2_x2_4_sig
* NET 706 = no4_x1_3_sig
* NET 707 = aux38
* NET 708 = o3_x2_4_sig
* NET 711 = not_cuh[1]
* NET 716 = cum_1_ins.sff_s
* NET 718 = cum_1_ins.y
* NET 719 = cum_1_ins.u
* NET 722 = cum_1_ins.sff_m
* NET 724 = cum_1_ins.ckr
* NET 725 = cum_1_ins.nckr
* NET 728 = not_cum[0]
* NET 730 = not_cuh[3]
* NET 731 = not_aux1
* NET 736 = not_cum[3]
* NET 740 = oa22_x2_17_sig
* NET 741 = on12_x1_7_sig
* NET 746 = xr2_x1_3_sig
* NET 750 = not_cdm[3]
* NET 758 = na3_x1_8_sig
* NET 759 = not_aux38
* NET 761 = not_cum[1]
* NET 762 = mbk_buf_not_cum[3]
* NET 766 = rtlalc_10_0_ins.ckr
* NET 767 = rtlalc_10_0_ins.nckr
* NET 768 = rtlalc_10_0_ins.sff_s
* NET 770 = rtlalc_10_0_ins.sff_m
* NET 771 = rtlalc_10_0_ins.y
* NET 774 = rtlalc_10_0_ins.u
* NET 778 = na2_x1_7_sig
* NET 779 = na4_x1_4_sig
* NET 780 = na2_x1_8_sig
* NET 785 = ao2o22_x2_5_sig
* NET 788 = not_aux43
* NET 793 = oa22_x2_6_sig
* NET 794 = on12_x1_2_sig
* NET 798 = a2_x2_3_sig
* NET 801 = cuh[0]
* NET 802 = cuh_0_ins.ckr
* NET 803 = cuh_0_ins.nckr
* NET 804 = cuh_0_ins.sff_m
* NET 806 = cuh_0_ins.sff_s
* NET 807 = cuh_0_ins.y
* NET 809 = noa22_x1_8_sig
* NET 812 = cuh_0_ins.u
* NET 818 = na3_x1_12_sig
* NET 819 = maquina
* NET 820 = nao22_x1_3_sig
* NET 823 = na3_x1_13_sig
* NET 824 = nao22_x1_4_sig
* NET 828 = o2_x2_6_sig
* NET 829 = not_aux68
* NET 830 = not_aux119
* NET 833 = not_cum[2]
* NET 834 = on12_x1_6_sig
* NET 839 = dh[0]
* NET 841 = uh[2]
* NET 843 = rtlalc_10[0]
* NET 845 = uh[1]
* NET 846 = uh[0]
* NET 848 = rtlalc_10[3]
* NET 850 = rtlalc_10_3_ins.sff_m
* NET 851 = rtlalc_10_3_ins.y
* NET 852 = rtlalc_10_3_ins.sff_s
* NET 854 = rtlalc_10_3_ins.u
* NET 855 = rtlalc_10_3_ins.ckr
* NET 856 = rtlalc_10_3_ins.nckr
* NET 860 = a2_x2_4_sig
* NET 861 = no3_x1_sig
* NET 862 = aux49
* NET 864 = rtlalc_10[2]
* NET 866 = rtlalc_10_2_ins.sff_s
* NET 867 = rtlalc_10_2_ins.y
* NET 868 = rtlalc_10_2_ins.u
* NET 870 = rtlalc_10_2_ins.sff_m
* NET 872 = rtlalc_10_2_ins.ckr
* NET 873 = rtlalc_10_2_ins.nckr
* NET 874 = a3_x2_sig
* NET 875 = nao22_x1_2_sig
* NET 878 = not_cuh[0]
* NET 880 = inv_x2_6_sig
* NET 881 = not_aux42
* NET 883 = oa22_x2_10_sig
* NET 884 = noa22_x1_12_sig
* NET 887 = oa22_x2_9_sig
* NET 889 = ao2o22_x2_8_sig
* NET 890 = mbk_buf_not_cuh[3]
* NET 893 = cuh[3]
* NET 895 = cuh_3_ins.sff_s
* NET 897 = cuh_3_ins.y
* NET 898 = noa22_x1_11_sig
* NET 899 = cuh_3_ins.u
* NET 900 = cuh_3_ins.sff_m
* NET 902 = cuh_3_ins.ckr
* NET 903 = cuh_3_ins.nckr
* NET 907 = nao2o22_x1_sig
* NET 908 = not_aux113
* NET 909 = a3_x2_5_sig
* NET 912 = aux69
* NET 915 = not_maquina
* NET 919 = mdh_1_ins.sff_m
* NET 920 = mdh_1_ins.sff_s
* NET 921 = mdh_1_ins.y
* NET 923 = mdh_1_ins.u
* NET 924 = mdh_1_ins.ckr
* NET 925 = mdh_1_ins.nckr
* NET 949 = dm[3]
* NET 950 = rtlalc_11[3]
* NET 952 = rtlalc_11_3_ins.y
* NET 954 = rtlalc_11_3_ins.sff_m
* NET 955 = rtlalc_11_3_ins.sff_s
* NET 957 = rtlalc_11_3_ins.u
* NET 959 = rtlalc_11_3_ins.ckr
* NET 962 = ao2o22_x2_12_sig
* NET 963 = rtlalc_11_3_ins.nckr
* NET 965 = cdm[3]
* NET 969 = rtlalc_10[1]
* NET 971 = rtlalc_10_1_ins.y
* NET 972 = rtlalc_10_1_ins.sff_s
* NET 975 = rtlalc_10_1_ins.u
* NET 977 = rtlalc_10_1_ins.sff_m
* NET 978 = rtlalc_10_1_ins.ckr
* NET 980 = rtlalc_9[0]
* NET 981 = rtlalc_10_1_ins.nckr
* NET 985 = rtlalc_9_0_ins.sff_s
* NET 986 = rtlalc_9_0_ins.y
* NET 988 = rtlalc_9_0_ins.ckr
* NET 989 = rtlalc_9_0_ins.u
* NET 991 = rtlalc_9_0_ins.sff_m
* NET 992 = rtlalc_9_0_ins.nckr
* NET 993 = ao2o22_x2_6_sig
* NET 995 = cuh[1]
* NET 1001 = ao2o22_x2_7_sig
* NET 1003 = cuh[2]
* NET 1007 = cdm[1]
* NET 1012 = ao2o22_x2_sig
* NET 1015 = cdh[0]
* NET 1018 = cum[1]
* NET 1024 = cum_2_ins.sff_s
* NET 1026 = cum_2_ins.y
* NET 1027 = oa22_x2_16_sig
* NET 1029 = cum_2_ins.sff_m
* NET 1031 = cum_2_ins.nckr
* NET 1032 = cum_2_ins.u
* NET 1033 = cum_2_ins.ckr
* NET 1042 = oa2a2a23_x2_sig
* NET 1043 = no2_x1_9_sig
* NET 1044 = aux77
* NET 1047 = no2_x1_7_sig
* NET 1050 = not_aux77
* NET 1052 = nao2o22_x1_2_sig
* NET 1057 = o4_x2_4_sig
* NET 1061 = dm[2]
* NET 1064 = rtlalc_11[2]
* NET 1066 = rtlalc_11_2_ins.sff_s
* NET 1067 = rtlalc_11_2_ins.y
* NET 1070 = rtlalc_11_2_ins.sff_m
* NET 1071 = rtlalc_11_2_ins.ckr
* NET 1072 = rtlalc_11_2_ins.nckr
* NET 1073 = rtlalc_11_2_ins.u
* NET 1075 = rtlalc_12[1]
* NET 1076 = rtlalc_12_1_ins.sff_s
* NET 1077 = ao2o22_x2_14_sig
* NET 1078 = rtlalc_12_1_ins.y
* NET 1079 = rtlalc_12_1_ins.u
* NET 1080 = rtlalc_12_1_ins.sff_m
* NET 1083 = rtlalc_12_1_ins.ckr
* NET 1084 = rtlalc_12_1_ins.nckr
* NET 1085 = ao2o22_x2_11_sig
* NET 1086 = cdm[2]
* NET 1092 = mdh_3_ins.sff_s
* NET 1093 = mdh_3_ins.y
* NET 1095 = mdh_3_ins.sff_m
* NET 1097 = mdh_3_ins.ckr
* NET 1098 = mdh_3_ins.nckr
* NET 1099 = mdh_3_ins.u
* NET 1100 = oa2ao222_x2_2_sig
* NET 1104 = aux122
* NET 1110 = xr2_x1_4_sig
* NET 1114 = mbk_buf_aux74
* NET 1115 = mdh[2]
* NET 1117 = mdh_2_ins.y
* NET 1118 = mdh_2_ins.sff_s
* NET 1119 = mdh_2_ins.sff_m
* NET 1122 = oa2a22_x2_sig
* NET 1123 = mdh_2_ins.u
* NET 1124 = mdh_2_ins.ckr
* NET 1125 = mdh_2_ins.nckr
* NET 1127 = na2_x1_17_sig
* NET 1128 = no2_x1_8_sig
* NET 1129 = na4_x1_6_sig
* NET 1133 = no3_x1_3_sig
* NET 1134 = na2_x1_19_sig
* NET 1157 = dm[1]
* NET 1160 = rtlalc_11_0_ins.y
* NET 1162 = rtlalc_11_0_ins.sff_s
* NET 1163 = rtlalc_11_0_ins.ckr
* NET 1164 = rtlalc_11_0_ins.u
* NET 1165 = rtlalc_11_0_ins.sff_m
* NET 1167 = ao2o22_x2_9_sig
* NET 1168 = rtlalc_11_0_ins.nckr
* NET 1169 = cdm[0]
* NET 1173 = cum[2]
* NET 1177 = not_mdh[2]
* NET 1178 = inv_x2_9_sig
* NET 1185 = no4_x1_6_sig
* NET 1187 = a2_x2_9_sig
* NET 1188 = xr2_x1_5_sig
* NET 1190 = rtlalc_11[1]
* NET 1192 = rtlalc_11_1_ins.sff_s
* NET 1193 = ao2o22_x2_10_sig
* NET 1194 = rtlalc_11_1_ins.y
* NET 1196 = rtlalc_11_1_ins.sff_m
* NET 1198 = rtlalc_11_1_ins.nckr
* NET 1199 = rtlalc_11_1_ins.ckr
* NET 1200 = rtlalc_11_1_ins.u
* NET 1201 = mdh[3]
* NET 1202 = a2_x2_8_sig
* NET 1204 = not_muh[0]
* NET 1206 = aux79
* NET 1207 = aux74
* NET 1208 = inv_x2_sig
* NET 1213 = mdh_0_ins.sff_s
* NET 1214 = mdh_0_ins.y
* NET 1216 = mdh_0_ins.sff_m
* NET 1218 = mdh_0_ins.u
* NET 1219 = mdh_0_ins.nckr
* NET 1220 = mdh_0_ins.ckr
* NET 1221 = oa22_x2_18_sig
* NET 1224 = a3_x2_7_sig
* NET 1225 = aux70
* NET 1226 = inv_x2_8_sig
* NET 1228 = dm[0]
* NET 1229 = rtlalc_11[0]
* NET 1234 = rtlalc_12_3_ins.u
* NET 1235 = rtlalc_12_3_ins.ckr
* NET 1238 = rtlalc_12_3_ins.nckr
* NET 1239 = cum[0]
* NET 1241 = oa2a22_x2_5_sig
* NET 1243 = not_ctrl
* NET 1244 = ctrl
* NET 1245 = cum[3]
* NET 1257 = nao22_x1_7_sig
* NET 1259 = mdm_0_ins.ckr
* NET 1260 = mdm_0_ins.u
* NET 1264 = mdm_0_ins.nckr
* NET 1265 = aux123
* NET 1267 = not_aux87
* NET 1271 = na4_x1_sig
* NET 1276 = no2_x1_6_sig
* NET 1281 = no3_x1_2_sig
* NET 1282 = mbk_buf_not_aux74
* NET 1286 = nao22_x1_5_sig
* NET 1288 = na2_x1_18_sig
* NET 1293 = o4_x2_5_sig
* NET 1296 = rtlalc_12_3_ins.sff_s
* NET 1297 = rtlalc_12_3_ins.y
* NET 1298 = rtlalc_12_3_ins.sff_m
* NET 1308 = mdm[0]
* NET 1310 = nxr2_x1_3_sig
* NET 1311 = mdm_0_ins.sff_s
* NET 1313 = mdm_0_ins.y
* NET 1314 = mdm_0_ins.sff_m
* NET 1325 = mdh[1]
* NET 1326 = mdh[0]
* NET 1333 = not_aux74
* NET 1337 = na2_x1_16_sig
* NET 1338 = a3_x2_8_sig
* NET 1344 = rtlalc_12[3]
* NET 1345 = um[3]
* NET 1349 = rtlalc_12[0]
* NET 1350 = rtlalc_12_0_ins.y
* NET 1351 = rtlalc_12_0_ins.sff_s
* NET 1353 = ao2o22_x2_13_sig
* NET 1354 = rtlalc_12_0_ins.u
* NET 1356 = rtlalc_12_0_ins.sff_m
* NET 1357 = rtlalc_12_0_ins.ckr
* NET 1359 = rtlalc_12[2]
* NET 1360 = rtlalc_12_0_ins.nckr
* NET 1361 = rtlalc_12_2_ins.y
* NET 1363 = rtlalc_12_2_ins.sff_s
* NET 1365 = ao2o22_x2_15_sig
* NET 1366 = rtlalc_12_2_ins.u
* NET 1368 = rtlalc_12_2_ins.sff_m
* NET 1369 = rtlalc_12_2_ins.ckr
* NET 1370 = o3_x2_12_sig
* NET 1371 = rtlalc_12_2_ins.nckr
* NET 1375 = na2_x1_23_sig
* NET 1376 = not_aux98
* NET 1380 = aux98
* NET 1382 = on12_x1_8_sig
* NET 1384 = nao2o22_x1_4_sig
* NET 1387 = mdm_2_ins.y
* NET 1388 = mdm_2_ins.sff_s
* NET 1390 = oa22_x2_20_sig
* NET 1391 = mdm_2_ins.u
* NET 1394 = mdm_2_ins.sff_m
* NET 1395 = mdm_2_ins.ckr
* NET 1396 = mdm_2_ins.nckr
* NET 1400 = no4_x1_7_sig
* NET 1403 = no2_x1_13_sig
* NET 1405 = na4_x1_5_sig
* NET 1406 = o2_x2_10_sig
* NET 1409 = not_aux120
* NET 1410 = not_muh[3]
* NET 1414 = not_aux76
* NET 1415 = no2_x1_5_sig
* NET 1417 = not_aux75
* NET 1421 = muh_3_ins.sff_s
* NET 1422 = muh_3_ins.y
* NET 1424 = muh_3_ins.sff_m
* NET 1425 = oa2a22_x2_3_sig
* NET 1426 = muh_3_ins.u
* NET 1428 = muh_3_ins.nckr
* NET 1429 = muh_3_ins.ckr
* NET 1442 = aux124
* NET 1453 = no4_x1_8_sig
* NET 1468 = inv_x2_11_sig
* NET 1474 = um[2]
* NET 1475 = mdm_3_ins.sff_s
* NET 1476 = mdm_3_ins.sff_m
* NET 1477 = mdm_3_ins.y
* NET 1479 = mdm_3_ins.ckr
* NET 1480 = mdm_3_ins.u
* NET 1484 = mdm_3_ins.nckr
* NET 1485 = aux108
* NET 1487 = oa2a22_x2_4_sig
* NET 1489 = no2_x1_14_sig
* NET 1495 = xr2_x1_8_sig
* NET 1498 = aux105
* NET 1500 = not_aux105
* NET 1501 = an12_x1_4_sig
* NET 1502 = not_aux130
* NET 1504 = not_aux127
* NET 1506 = o2_x2_11_sig
* NET 1508 = not_aux106
* NET 1510 = mdm_1_ins.sff_s
* NET 1513 = mdm_1_ins.ckr
* NET 1514 = mdm_1_ins.u
* NET 1515 = mdm_1_ins.sff_m
* NET 1517 = mdm_1_ins.y
* NET 1518 = mdm_1_ins.nckr
* NET 1519 = nao2o22_x1_3_sig
* NET 1520 = na3_x1_sig
* NET 1523 = no2_x1_12_sig
* NET 1524 = na2_x1_21_sig
* NET 1528 = na4_x1_7_sig
* NET 1530 = na2_x1_22_sig
* NET 1535 = nxr2_x1_2_sig
* NET 1536 = not_aux78
* NET 1538 = nao22_x1_6_sig
* NET 1542 = muh_2_ins.sff_s
* NET 1543 = muh[2]
* NET 1544 = muh_2_ins.sff_m
* NET 1545 = muh_2_ins.ckr
* NET 1547 = muh_2_ins.y
* NET 1548 = muh_2_ins.nckr
* NET 1549 = muh_2_ins.u
* NET 1550 = oa2ao222_x2_4_sig
* NET 1552 = mum_1_ins.sff_s
* NET 1554 = mum_1_ins.y
* NET 1556 = mum_1_ins.sff_m
* NET 1558 = mum_1_ins.nckr
* NET 1559 = mum_1_ins.u
* NET 1560 = mum_1_ins.ckr
* NET 1562 = oa22_x2_21_sig
* NET 1564 = a3_x2_9_sig
* NET 1567 = o2_x2_12_sig
* NET 1569 = mdm[3]
* NET 1570 = not_mum[0]
* NET 1574 = not_mdm[0]
* NET 1575 = not_mum[3]
* NET 1578 = not_aux109
* NET 1579 = not_aux89
* NET 1581 = mdm[2]
* NET 1582 = not_aux73
* NET 1585 = not_mdm[1]
* NET 1586 = muh[3]
* NET 1587 = na2_x1_20_sig
* NET 1590 = no3_x1_4_sig
* NET 1594 = not_aux103
* NET 1596 = o2_x2_9_sig
* NET 1598 = noa22_x1_20_sig
* NET 1600 = a2_x2_12_sig
* NET 1601 = not_mdm[2]
* NET 1602 = not_aux96
* NET 1605 = not_mdh[0]
* NET 1607 = um[1]
* NET 1629 = mum_0_ins.y
* NET 1630 = mum_0_ins.sff_s
* NET 1633 = mum_0_ins.u
* NET 1635 = mum_0_ins.sff_m
* NET 1639 = mum_0_ins.nckr
* NET 1640 = mum_0_ins.ckr
* NET 1641 = aux111
* NET 1646 = aux110
* NET 1650 = mum[0]
* NET 1654 = aux73
* NET 1657 = mbk_buf_aux73
* NET 1664 = xr2_x1_6_sig
* NET 1670 = no2_x1_10_sig
* NET 1672 = not_aux90
* NET 1673 = a2_x2_10_sig
* NET 1677 = mbk_buf_not_mum[3]
* NET 1681 = muh_0_ins.y
* NET 1684 = muh_0_ins.sff_m
* NET 1686 = muh_0_ins.sff_s
* NET 1687 = oa2a22_x2_2_sig
* NET 1688 = muh_0_ins.u
* NET 1689 = muh_0_ins.ckr
* NET 1690 = muh_0_ins.nckr
* NET 1695 = a2_x2_sig
* NET 1696 = not_aux102
* NET 1701 = na2_x1_sig
* NET 1707 = a2_x2_11_sig
* NET 1708 = rst
* NET 1709 = not_aux121
* NET 1710 = mdm[1]
* NET 1715 = not_aux125
* NET 1716 = o3_x2_11_sig
* NET 1719 = o2_x2_8_sig
* NET 1722 = oa22_x2_19_sig
* NET 1726 = o2_x2_7_sig
* NET 1727 = vss
* NET 1728 = um[0]
* NET 1730 = mum_2_ins.sff_s
* NET 1731 = mum_2_ins.y
* NET 1733 = mum_2_ins.u
* NET 1735 = mum_2_ins.sff_m
* NET 1736 = oa22_x2_22_sig
* NET 1737 = mum_2_ins.nckr
* NET 1738 = mum_2_ins.ckr
* NET 1739 = mx2_x2_sig
* NET 1742 = a3_x2_10_sig
* NET 1746 = mum_3_ins.sff_s
* NET 1747 = mum_3_ins.y
* NET 1748 = mum_3_ins.ckr
* NET 1749 = mum_3_ins.u
* NET 1751 = mum_3_ins.sff_m
* NET 1752 = mum[3]
* NET 1753 = mum_3_ins.nckr
* NET 1757 = xr2_x1_9_sig
* NET 1758 = not_rst
* NET 1759 = oa22_x2_23_sig
* NET 1762 = na3_x1_15_sig
* NET 1764 = nao22_x1_8_sig
* NET 1765 = a3_x2_11_sig
* NET 1766 = inv_x2_12_sig
* NET 1767 = aux112
* NET 1769 = mbk_buf_mum[0]
* NET 1770 = na2_x1_24_sig
* NET 1771 = mum[1]
* NET 1772 = mum[2]
* NET 1776 = not_muh[2]
* NET 1778 = not_aux91
* NET 1780 = not_aux97
* NET 1781 = a2_x2_13_sig
* NET 1783 = not_mum[2]
* NET 1784 = no2_x1_11_sig
* NET 1785 = not_mum[1]
* NET 1786 = muh[0]
* NET 1790 = not_aux93
* NET 1791 = o3_x2_10_sig
* NET 1792 = not_muh[1]
* NET 1793 = na3_x1_14_sig
* NET 1795 = noa22_x1_18_sig
* NET 1796 = noa22_x1_19_sig
* NET 1797 = xr2_x1_7_sig
* NET 1801 = not_aux129
* NET 1802 = inv_x2_10_sig
* NET 1804 = muh_1_ins.sff_s
* NET 1805 = muh_1_ins.y
* NET 1807 = muh_1_ins.sff_m
* NET 1808 = muh[1]
* NET 1809 = oa2ao222_x2_3_sig
* NET 1810 = clk
* NET 1812 = muh_1_ins.u
* NET 1813 = muh_1_ins.ckr
* NET 1814 = vdd
* NET 1815 = muh_1_ins.nckr
Mtr_03624 1814 1791 1794 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03623 1795 1793 1794 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03622 1794 1792 1795 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03621 1802 1801 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03620 1809 1798 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03619 1800 1795 1799 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03618 1800 1802 1814 1814 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03617 1814 1808 1800 1814 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03616 1799 1796 1798 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03615 1798 1797 1800 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03614 1787 1786 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03613 1814 1808 1788 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03612 1797 1787 1789 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03611 1789 1808 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03610 1789 1788 1797 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03609 1814 1786 1789 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03608 1803 1808 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03607 1804 1813 1803 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03606 1805 1815 1804 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03605 1807 1815 1806 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03604 1806 1805 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03603 1811 1813 1807 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03602 1815 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03601 1814 1815 1813 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03600 1812 1809 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03599 1814 1812 1811 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03598 1814 1804 1808 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03597 1808 1804 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03596 1805 1807 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03595 1779 1778 1784 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03594 1814 1780 1779 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03593 1814 1778 1774 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03592 1774 1772 1773 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03591 1773 1771 1775 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03590 1790 1775 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03589 1814 1785 1793 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03588 1793 1783 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03587 1793 1784 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03586 1780 1777 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03585 1814 1776 1777 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03584 1777 1786 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03583 1781 1782 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03582 1814 1792 1782 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03581 1782 1780 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03580 1770 1769 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03579 1814 1783 1770 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03578 1814 1761 1759 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03577 1760 1765 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03576 1760 1764 1761 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03575 1761 1771 1760 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03574 1814 1770 1768 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03573 1765 1768 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03572 1814 1767 1768 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03571 1768 1785 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03570 1814 1762 1764 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03569 1763 1772 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03568 1764 1766 1763 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03567 1766 1767 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03566 1754 1752 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03565 1814 1769 1755 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03564 1757 1754 1756 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03563 1756 1769 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03562 1756 1755 1757 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03561 1814 1752 1756 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03560 1814 1772 1762 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03559 1762 1757 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03558 1762 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03557 1745 1752 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03556 1746 1748 1745 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03555 1747 1753 1746 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03554 1751 1753 1744 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03553 1744 1747 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03552 1750 1748 1751 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03551 1753 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03550 1814 1753 1748 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03549 1749 1759 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03548 1814 1749 1750 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03547 1814 1746 1752 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03546 1752 1746 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03545 1747 1751 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03544 1814 1785 1743 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03543 1742 1743 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03542 1814 1758 1743 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03541 1743 1772 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03540 1729 1772 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03539 1730 1738 1729 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03538 1731 1737 1730 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03537 1735 1737 1734 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03536 1734 1731 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03535 1732 1738 1735 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03534 1737 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03533 1814 1737 1738 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03532 1733 1736 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03531 1814 1733 1732 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03530 1814 1730 1772 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03529 1772 1730 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03528 1731 1735 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03527 1814 1741 1736 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03526 1740 1742 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03525 1740 1739 1741 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03524 1741 1771 1740 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03523 1814 1758 1801 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03522 1625 1790 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03521 1801 1710 1625 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03520 1814 1716 1626 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03519 1796 1722 1626 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03518 1626 1715 1796 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03517 1707 1704 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03516 1814 1792 1704 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03515 1704 1790 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03514 1814 1721 1722 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03513 1627 1726 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03512 1627 1719 1721 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03511 1721 1776 1627 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03510 1814 1708 1624 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03509 1624 1709 1623 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03508 1623 1707 1711 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03507 1716 1711 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03506 1792 1808 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03505 1814 1772 1622 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03504 1622 1701 1621 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03503 1621 1695 1697 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03502 1696 1697 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03501 1628 1771 1724 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03500 1814 1772 1628 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03499 1726 1724 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03498 1695 1693 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03497 1814 1776 1693 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03496 1693 1778 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03495 1701 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03494 1814 1785 1701 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03493 1657 1655 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03492 1814 1654 1655 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03491 1785 1771 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03490 1783 1772 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03489 1658 1786 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03488 1814 1657 1660 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03487 1664 1658 1614 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03486 1614 1657 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03485 1614 1660 1664 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03484 1814 1786 1614 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03483 1617 1677 1767 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03482 1814 1708 1617 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03481 1618 1786 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03480 1686 1689 1618 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03479 1681 1690 1686 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03478 1684 1690 1620 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03477 1620 1681 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03476 1619 1689 1684 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03475 1690 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03474 1814 1690 1689 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03473 1688 1687 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03472 1814 1688 1619 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03471 1814 1686 1786 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03470 1786 1686 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03469 1681 1684 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03468 1673 1674 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03467 1814 1758 1674 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03466 1674 1672 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03465 1615 1664 1665 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03464 1615 1670 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03463 1814 1786 1615 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03462 1665 1673 1615 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03461 1687 1665 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03460 1616 1672 1670 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03459 1814 1708 1616 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03458 1814 1644 1739 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03457 1612 1646 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03456 1649 1772 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03455 1611 1772 1644 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03454 1644 1649 1612 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03453 1814 1641 1611 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03452 1613 1769 1646 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03451 1814 1708 1613 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03450 1769 1651 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03449 1814 1650 1651 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03448 1608 1650 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03447 1630 1640 1608 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03446 1629 1639 1630 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03445 1635 1639 1610 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03444 1610 1629 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03443 1609 1640 1635 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03442 1639 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03441 1814 1639 1640 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03440 1633 1646 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03439 1814 1633 1609 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03438 1814 1630 1650 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03437 1650 1630 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03436 1629 1635 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03435 1604 1601 1603 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03434 1814 1602 1604 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03433 1719 1603 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03432 1591 1709 1592 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03431 1814 1696 1591 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03430 1596 1592 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03429 1715 1606 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03428 1814 1605 1606 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03427 1606 1808 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03426 1814 1596 1597 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03425 1598 1776 1597 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03424 1597 1600 1598 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03423 1600 1599 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03422 1814 1715 1599 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03421 1599 1602 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03420 1585 1710 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03419 1587 1586 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03418 1814 1585 1587 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03417 1593 1776 1595 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03416 1814 1808 1593 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03415 1594 1595 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03414 1814 1587 1589 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03413 1588 1781 1590 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03412 1589 1696 1588 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03411 1584 1582 1583 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03410 1814 1601 1584 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03409 1778 1583 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03408 1578 1579 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03407 1814 1710 1578 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03406 1814 1783 1580 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03405 1579 1580 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03404 1814 1581 1580 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03403 1580 1785 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03402 1672 1577 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03401 1814 1585 1577 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03400 1577 1579 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03399 1601 1581 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03398 1582 1654 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03397 1814 1567 1565 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03396 1564 1565 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03395 1814 1641 1565 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03394 1565 1785 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03393 1677 1576 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03392 1814 1575 1576 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03391 1814 1575 1573 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03390 1572 1569 1571 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03389 1571 1574 1654 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03388 1573 1570 1572 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03387 1570 1650 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03386 1566 1677 1568 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03385 1814 1772 1566 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03384 1567 1568 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03383 1575 1752 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03382 1814 1561 1562 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03381 1563 1564 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03380 1563 1771 1561 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03379 1561 1646 1563 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03378 1553 1771 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03377 1552 1560 1553 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03376 1554 1558 1552 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03375 1556 1558 1555 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03374 1555 1554 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03373 1557 1560 1556 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03372 1558 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03371 1814 1558 1560 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03370 1559 1562 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03369 1814 1559 1557 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03368 1814 1552 1771 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03367 1771 1552 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03366 1554 1556 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03365 1814 1594 1538 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03364 1462 1792 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03363 1538 1535 1462 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03362 1814 1531 1461 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03361 1461 1532 1535 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03360 1461 1543 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03359 1535 1786 1461 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03358 1814 1543 1532 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03357 1531 1786 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03356 1468 1801 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03355 1550 1539 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03354 1465 1598 1464 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03353 1465 1468 1814 1814 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03352 1814 1543 1465 1814 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03351 1464 1590 1539 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03350 1539 1538 1465 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03349 1469 1543 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03348 1542 1545 1469 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03347 1547 1548 1542 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03346 1544 1548 1471 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03345 1471 1547 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03344 1472 1545 1544 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03343 1548 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03342 1814 1548 1545 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03341 1549 1550 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03340 1814 1549 1472 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03339 1814 1542 1543 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03338 1543 1542 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03337 1547 1544 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03336 1814 1792 1520 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03335 1520 1585 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03334 1520 1776 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03333 1814 1785 1528 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03332 1528 1523 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03331 1814 1524 1528 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03330 1528 1783 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03329 1460 1710 1523 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03328 1814 1530 1460 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03327 1530 1594 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03326 1814 1536 1530 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03325 1524 1808 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03324 1814 1776 1524 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03323 1519 1501 1448 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03322 1448 1506 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03321 1447 1585 1519 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03320 1814 1502 1447 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03319 1449 1504 1503 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03318 1814 1508 1449 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03317 1506 1503 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03316 1497 1581 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03315 1814 1497 1445 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03314 1445 1569 1501 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03313 1814 1581 1450 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03312 1451 1585 1452 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03311 1452 1508 1453 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03310 1450 1771 1451 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03309 1454 1710 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03308 1510 1513 1454 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03307 1517 1518 1510 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03306 1515 1518 1457 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03305 1457 1517 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03304 1456 1513 1515 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03303 1518 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03302 1814 1518 1513 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03301 1514 1519 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03300 1814 1514 1456 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03299 1814 1510 1710 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03298 1710 1510 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03297 1517 1515 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03296 1446 1500 1499 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03295 1814 1708 1446 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03294 1508 1499 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03293 1437 1570 1641 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03292 1814 1708 1437 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03291 1500 1498 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03290 1441 1570 1442 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03289 1814 1677 1441 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03288 1814 1574 1443 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03287 1444 1570 1498 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03286 1443 1677 1444 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03285 1438 1495 1486 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03284 1438 1485 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03283 1814 1578 1438 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03282 1486 1489 1438 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03281 1487 1486 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03280 1435 1578 1489 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03279 1814 1708 1435 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03278 1491 1569 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03277 1814 1498 1492 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03276 1495 1491 1440 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03275 1440 1498 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03274 1440 1492 1495 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03273 1814 1569 1440 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03272 1430 1569 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03271 1475 1479 1430 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03270 1477 1484 1475 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03269 1476 1484 1433 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03268 1433 1477 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03267 1432 1479 1476 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03266 1484 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03265 1814 1484 1479 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03264 1480 1487 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03263 1814 1480 1432 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03262 1814 1475 1569 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03261 1569 1475 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03260 1477 1476 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03259 1416 1414 1415 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03258 1814 1409 1416 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03257 1814 1708 1411 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03256 1411 1710 1413 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03255 1413 1410 1412 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03254 1791 1412 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03253 1776 1543 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03252 1418 1417 1419 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03251 1814 1601 1418 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03250 1414 1419 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03249 1407 1414 1408 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03248 1814 1709 1407 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03247 1406 1408 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03246 1420 1586 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03245 1421 1429 1420 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03244 1422 1428 1421 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03243 1424 1428 1423 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03242 1423 1422 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03241 1427 1429 1424 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03240 1428 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03239 1814 1428 1429 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03238 1426 1425 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03237 1814 1426 1427 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03236 1814 1421 1586 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03235 1586 1421 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03234 1422 1424 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03233 1814 1415 1405 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03232 1405 1785 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03231 1814 1783 1405 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03230 1405 1776 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03229 1404 1410 1403 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03228 1814 1708 1404 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03227 1814 1771 1397 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03226 1398 1776 1399 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03225 1399 1792 1400 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03224 1397 1406 1398 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03223 1401 1403 1402 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03222 1401 1400 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03221 1814 1783 1401 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03220 1402 1528 1401 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03219 1425 1402 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03218 1814 1485 1382 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03217 1382 1379 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03216 1814 1504 1379 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03215 1384 1601 1383 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03214 1383 1382 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03213 1381 1601 1384 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03212 1814 1502 1381 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03211 1389 1581 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03210 1388 1395 1389 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03209 1387 1396 1388 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03208 1394 1396 1393 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03207 1393 1387 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03206 1392 1395 1394 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03205 1396 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03204 1814 1396 1395 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03203 1391 1390 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03202 1814 1391 1392 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03201 1814 1388 1581 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03200 1581 1388 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03199 1387 1394 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03198 1814 1386 1390 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03197 1385 1384 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03196 1385 1453 1386 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03195 1386 1783 1385 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03194 1380 1785 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03193 1814 1783 1380 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03192 1375 1376 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03191 1814 1758 1375 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03190 1814 1758 1502 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03189 1378 1500 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03188 1502 1380 1378 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03187 1352 1349 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03186 1351 1357 1352 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03185 1350 1360 1351 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03184 1356 1360 1358 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03183 1358 1350 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03182 1355 1357 1356 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03181 1360 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03180 1814 1360 1357 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03179 1354 1353 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03178 1814 1354 1355 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03177 1814 1351 1349 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03176 1349 1351 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03175 1350 1356 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03174 1814 1708 1372 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03173 1372 1376 1373 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03172 1373 1574 1374 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03171 1370 1374 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03170 1376 1380 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03169 1474 1347 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03168 1814 1359 1347 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03167 1728 1348 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03166 1814 1349 1348 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03165 1364 1359 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03164 1363 1369 1364 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03163 1361 1371 1363 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03162 1368 1371 1362 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03161 1362 1361 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03160 1367 1369 1368 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03159 1371 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03158 1814 1371 1369 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03157 1366 1365 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03156 1814 1366 1367 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03155 1814 1363 1359 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03154 1359 1363 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03153 1361 1368 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03152 1345 1346 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03151 1814 1344 1346 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03150 1485 1377 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03149 1814 1569 1377 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03148 1377 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03147 1814 1333 1334 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03146 1814 1334 1282 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03145 1282 1334 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03144 1814 1334 1282 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03143 1282 1334 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03142 1283 1282 1536 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03141 1814 1601 1283 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03140 1605 1326 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03139 1291 1601 1339 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03138 1292 1417 1291 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03137 1290 1325 1292 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03136 1814 1605 1290 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03135 1814 1339 1293 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03134 1294 1808 1341 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03133 1814 1326 1294 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03132 1409 1341 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03131 1288 1409 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03130 1814 1536 1288 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03129 1275 1771 1276 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03128 1814 1808 1275 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03127 1814 1405 1286 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03126 1284 1337 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03125 1286 1338 1284 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03124 1814 1281 1329 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03123 1338 1329 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03122 1814 1783 1329 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03121 1329 1276 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03120 1337 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03119 1814 1326 1337 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03118 1814 1282 1280 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03117 1279 1543 1281 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03116 1280 1601 1279 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03115 1265 1319 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03114 1814 1758 1319 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03113 1319 1267 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03112 1758 1708 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03111 1270 1520 1322 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03110 1268 1771 1270 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03109 1269 1772 1268 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03108 1814 1271 1269 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03107 1814 1322 1267 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03106 1814 1325 1271 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03105 1271 1326 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03104 1814 1581 1271 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03103 1271 1586 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03102 1814 1710 1262 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03101 1262 1772 1263 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03100 1263 1771 1317 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03099 1504 1317 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03098 1182 1308 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03097 1311 1259 1182 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03096 1313 1264 1311 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03095 1314 1264 1254 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03094 1254 1313 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03093 1258 1259 1314 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03092 1264 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03091 1814 1264 1259 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03090 1260 1257 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03089 1814 1260 1258 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03088 1814 1311 1308 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03087 1308 1311 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03086 1313 1314 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03085 1814 1306 1249 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03084 1249 1307 1310 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03083 1249 1442 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03082 1310 1308 1249 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03081 1814 1442 1307 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03080 1306 1308 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03079 1240 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03078 1237 1769 1300 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03077 1814 1244 1237 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03076 1300 1239 1240 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03075 1353 1300 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03074 1814 1370 1257 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03073 1252 1375 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03072 1257 1310 1252 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03071 1246 1245 1303 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03070 1246 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03069 1814 1752 1246 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03068 1303 1244 1246 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03067 1241 1303 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03066 1228 1295 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03065 1814 1229 1295 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03064 1158 1344 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03063 1296 1235 1158 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03062 1297 1238 1296 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03061 1298 1238 1231 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03060 1231 1297 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03059 1233 1235 1298 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03058 1238 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03057 1814 1238 1235 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03056 1234 1241 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03055 1814 1234 1233 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03054 1814 1296 1344 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03053 1344 1296 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03052 1297 1298 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03051 1212 1326 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03050 1213 1220 1212 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03049 1214 1219 1213 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03048 1216 1219 1217 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03047 1217 1214 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03046 1215 1220 1216 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03045 1219 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03044 1814 1219 1220 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03043 1218 1221 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03042 1814 1218 1215 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03041 1814 1213 1326 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03040 1326 1213 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03039 1214 1216 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03038 1226 1225 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03037 1814 1226 1227 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03036 1224 1227 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03035 1814 1758 1227 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03034 1227 1326 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03033 1210 1333 1211 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03032 1814 1708 1210 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03031 1417 1211 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03030 1814 1222 1221 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03029 1223 1224 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03028 1223 1286 1222 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03027 1222 1225 1223 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03026 1205 1582 1207 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03025 1814 1204 1205 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03024 1208 1206 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03023 1333 1207 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03022 1202 1203 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03021 1814 1204 1203 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03020 1203 1201 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03019 1204 1786 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03018 1814 1208 1209 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03017 1602 1209 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03016 1814 1325 1209 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03015 1209 1786 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03014 1191 1190 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03013 1192 1199 1191 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03012 1194 1198 1192 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03011 1196 1198 1197 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03010 1197 1194 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03009 1195 1199 1196 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03008 1198 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03007 1814 1198 1199 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03006 1200 1193 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03005 1814 1200 1195 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03004 1814 1192 1190 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03003 1190 1192 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03002 1194 1196 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03001 1184 1201 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03000 1814 1185 1186 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02999 1188 1184 1183 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02998 1183 1185 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02997 1183 1186 1188 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02996 1814 1201 1183 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02995 1187 1189 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02994 1814 1786 1189 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02993 1189 1188 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02992 1814 1569 1179 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02991 1180 1177 1181 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02990 1181 1178 1185 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02989 1179 1574 1180 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02988 1574 1308 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02987 1175 1244 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02986 1174 1173 1176 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02985 1814 1243 1174 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02984 1176 1772 1175 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02983 1365 1176 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02982 1170 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02981 1172 1308 1171 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02980 1814 1244 1172 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02979 1171 1169 1170 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02978 1167 1171 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02977 1178 1442 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02976 1159 1229 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02975 1162 1163 1159 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02974 1160 1168 1162 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02973 1165 1168 1161 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02972 1161 1160 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02971 1166 1163 1165 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02970 1168 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02969 1814 1168 1163 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02968 1164 1167 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02967 1814 1164 1166 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02966 1814 1162 1229 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02965 1229 1162 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02964 1160 1165 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02963 1157 1156 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02962 1814 1190 1156 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02961 1127 1808 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02960 1814 1206 1127 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02959 1046 1710 1128 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02958 1814 1288 1046 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02957 1814 1543 1054 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02956 1055 1772 1133 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02955 1054 1771 1055 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02954 1814 1128 1129 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02953 1129 1133 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02952 1814 1127 1129 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02951 1129 1134 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02950 1134 1326 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02949 1814 1808 1134 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02948 1410 1586 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02947 1814 1177 1206 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02946 1206 1090 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02945 1814 1201 1090 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02944 1114 1113 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02943 1814 1207 1113 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02942 1108 1115 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02941 1814 1114 1112 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02940 1110 1108 1025 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02939 1025 1114 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02938 1025 1112 1110 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02937 1814 1115 1025 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02936 1177 1115 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02935 1034 1115 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02934 1118 1124 1034 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02933 1117 1125 1118 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02932 1119 1125 1037 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02931 1037 1117 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02930 1038 1124 1119 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02929 1125 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02928 1814 1125 1124 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02927 1123 1122 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02926 1814 1123 1038 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02925 1814 1118 1115 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02924 1115 1118 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02923 1117 1119 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02922 1014 1267 1104 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02921 1814 1708 1014 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02920 1100 1103 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02919 1011 1202 1006 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02918 1011 1265 1814 1814 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02917 1814 1201 1011 1814 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02916 1006 1187 1103 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02915 1103 1104 1011 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02914 994 1201 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02913 1092 1097 994 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02912 1093 1098 1092 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02911 1095 1098 1000 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02910 1000 1093 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02909 999 1097 1095 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02908 1098 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02907 1814 1098 1097 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02906 1099 1100 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02905 1814 1099 999 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02904 1814 1092 1201 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02903 1201 1092 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02902 1093 1095 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02901 1021 1110 1106 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02900 1021 1265 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02899 1814 1115 1021 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02898 1106 1104 1021 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02897 1122 1106 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02896 982 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02895 983 1581 1087 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02894 1814 1244 983 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02893 1087 1086 982 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02892 1085 1087 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02891 968 1075 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02890 1076 1083 968 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02889 1078 1084 1076 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02888 1080 1084 974 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02887 974 1078 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02886 973 1083 1080 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02885 1084 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02884 1814 1084 1083 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02883 1079 1077 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02882 1814 1079 973 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02881 1814 1076 1075 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02880 1075 1076 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02879 1078 1080 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02878 956 1064 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02877 1066 1071 956 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02876 1067 1072 1066 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02875 1070 1072 961 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02874 961 1067 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02873 960 1071 1070 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02872 1072 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02871 1814 1072 1071 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02870 1073 1085 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02869 1814 1073 960 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02868 1814 1066 1064 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02867 1064 1066 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02866 1067 1070 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02865 1607 1062 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02864 1814 1075 1062 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02863 1061 1063 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02862 1814 1064 1063 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02861 1040 1410 1225 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02860 1814 1710 1040 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02859 1041 1709 1043 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02858 1814 1050 1041 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02857 1052 1057 1053 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02856 1053 1293 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02855 1051 1050 1052 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02854 1814 1326 1051 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02853 1042 1049 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02852 1814 1326 1045 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02851 1045 1043 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02850 1045 1129 1048 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02849 1048 1044 1045 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02848 1049 1047 1048 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02847 1048 1052 1049 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02846 1059 1771 1058 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02845 1060 1543 1059 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02844 1056 1808 1060 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02843 1814 1772 1056 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02842 1814 1058 1057 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02841 1039 1410 1047 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02840 1814 1710 1039 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02839 1035 1710 1036 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02838 1814 1586 1035 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02837 1709 1036 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02836 1023 1173 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02835 1024 1033 1023 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02834 1026 1031 1024 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02833 1029 1031 1030 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02832 1030 1026 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02831 1028 1033 1029 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02830 1031 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02829 1814 1031 1033 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02828 1032 1027 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02827 1814 1032 1028 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02826 1814 1024 1173 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02825 1173 1024 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02824 1026 1029 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02823 1243 1244 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02822 1022 1244 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02821 1020 1018 1019 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02820 1814 1243 1020 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02819 1019 1771 1022 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02818 1077 1019 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02817 996 1244 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02816 998 995 997 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02815 1814 1243 998 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02814 997 1808 996 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02813 993 997 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02812 1009 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02811 1008 1710 1010 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02810 1814 1244 1008 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02809 1010 1007 1009 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02808 1193 1010 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02807 1005 1244 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02806 1002 1003 1004 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02805 1814 1243 1002 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02804 1004 1543 1005 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02803 1001 1004 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02802 1017 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02801 1013 1326 1016 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02800 1814 1244 1013 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02799 1016 1015 1017 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02798 1012 1016 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02797 970 969 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02796 972 978 970 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02795 971 981 972 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02794 977 981 979 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02793 979 971 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02792 976 978 977 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02791 981 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02790 1814 981 978 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02789 975 993 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02788 1814 975 976 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02787 1814 972 969 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02786 969 972 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02785 971 977 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02784 967 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02783 964 1569 966 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02782 1814 1244 964 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02781 966 965 967 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02780 962 966 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02779 984 980 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02778 985 988 984 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02777 986 992 985 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02776 991 992 987 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02775 987 986 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02774 990 988 991 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02773 992 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02772 1814 992 988 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02771 989 1012 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02770 1814 989 990 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02769 1814 985 980 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02768 980 985 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02767 986 991 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02766 951 950 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02765 955 959 951 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02764 952 963 955 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02763 954 963 953 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02762 953 952 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02761 958 959 954 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02760 963 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02759 1814 963 959 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02758 957 962 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02757 1814 957 958 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02756 1814 955 950 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02755 950 955 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02754 952 954 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02753 949 948 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02752 1814 950 948 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02751 836 1325 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02750 920 924 836 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02749 921 925 920 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02748 919 925 837 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02747 837 921 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02746 838 924 919 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02745 925 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02744 1814 925 924 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02743 923 1042 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02742 1814 923 838 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02741 1814 920 1325 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02740 1325 920 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02739 921 919 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02738 912 914 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02737 1814 1239 914 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02736 914 1018 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02735 916 1325 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02734 1814 916 832 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02733 832 1708 1044 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02732 1050 1044 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02731 1814 915 905 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02730 909 905 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02729 1814 1758 905 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02728 905 1173 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02727 880 908 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02726 816 893 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02725 895 902 816 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02724 897 903 895 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02723 900 903 817 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02722 817 897 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02721 822 902 900 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02720 903 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02719 1814 903 902 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02718 899 898 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02717 1814 899 822 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02716 1814 895 893 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02715 893 895 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02714 897 900 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02713 1814 911 1027 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02712 826 909 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02711 826 907 911 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02710 911 908 826 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02709 814 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02708 813 1586 891 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02707 1814 1244 813 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02706 891 893 814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02705 889 891 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02704 1814 880 799 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02703 884 893 799 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02702 799 881 884 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02701 796 878 879 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02700 1814 1173 796 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02699 881 879 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02698 1814 887 800 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02697 898 883 800 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02696 800 884 898 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02695 786 864 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02694 866 872 786 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02693 867 873 866 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02692 870 873 790 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02691 790 867 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02690 789 872 870 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02689 873 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02688 1814 873 872 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02687 868 1001 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02686 1814 868 789 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02685 1814 866 864 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02684 864 866 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02683 867 870 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02682 1814 885 887 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02681 808 1708 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02680 808 915 885 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02679 885 890 808 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02678 1814 877 883 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02677 792 881 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02676 792 874 877 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02675 877 875 792 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02674 775 848 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02673 852 855 775 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02672 851 856 852 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02671 850 856 776 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02670 776 851 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02669 777 855 850 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02668 856 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02667 1814 856 855 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02666 854 889 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02665 1814 854 777 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02664 1814 852 848 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02663 848 852 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02662 851 850 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02661 1814 860 875 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02660 782 862 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02659 875 861 782 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02658 860 859 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02657 1814 1086 859 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02656 859 995 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02655 845 847 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02654 1814 969 847 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02653 846 844 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02652 1814 843 844 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02651 841 842 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02650 1814 864 842 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02649 839 840 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02648 1814 980 840 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02647 915 819 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02646 763 762 827 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02645 1814 830 763 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02644 828 827 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02643 1814 1758 834 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02642 834 765 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02641 1814 912 765 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02640 907 833 835 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02639 835 834 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02638 831 829 907 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02637 1814 830 831 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02636 1814 1239 823 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02635 823 761 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02634 823 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02633 1814 818 820 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02632 821 819 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02631 820 829 821 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02630 1814 828 818 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02629 818 824 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02628 818 908 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02627 760 761 815 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02626 1814 1708 760 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02625 829 815 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02624 1814 823 824 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02623 825 1239 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02622 824 829 825 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02621 1814 878 758 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02620 758 833 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02619 758 759 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02618 1814 791 793 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02617 756 1708 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02616 756 915 791 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02615 791 878 756 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02614 1814 793 795 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02613 809 794 795 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02612 795 798 809 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02611 798 797 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02610 1814 908 797 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02609 797 758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02608 805 801 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02607 806 802 805 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02606 807 803 806 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02605 804 803 811 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02604 811 807 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02603 810 802 804 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02602 803 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02601 1814 803 802 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02600 812 809 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02599 1814 812 810 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02598 1814 806 801 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02597 801 806 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02596 807 804 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02595 778 1003 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02594 1814 750 778 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02593 755 915 787 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02592 1814 881 755 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02591 788 787 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02590 1814 778 783 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02589 781 779 861 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02588 783 780 781 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02587 754 1244 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02586 753 801 784 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02585 1814 1243 753 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02584 784 1786 754 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02583 785 784 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02582 780 1239 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02581 1814 1169 780 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02580 769 843 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02579 768 766 769 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02578 771 767 768 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02577 770 767 773 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02576 773 771 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02575 772 766 770 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02574 767 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02573 1814 767 766 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02572 774 785 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02571 1814 774 772 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02570 1814 768 843 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02569 843 768 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02568 771 770 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02567 750 965 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02566 1814 1245 736 1814 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02565 736 1245 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02564 762 737 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02563 1814 736 737 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02562 745 1245 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02561 1814 912 748 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02560 746 745 659 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02559 659 912 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02558 659 748 746 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02557 1814 1245 659 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02556 1814 739 740 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02555 658 1708 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02554 658 915 739 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02553 739 762 658 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02552 1814 746 741 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02551 741 744 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02550 1814 833 744 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02549 890 713 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02548 1814 730 713 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02547 1814 730 657 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02546 657 1018 656 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02545 656 736 733 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02544 731 733 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02543 711 995 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02542 652 1018 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02541 716 724 652 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02540 718 725 716 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02539 722 725 654 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02538 654 718 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02537 653 724 722 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02536 725 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02535 1814 725 724 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02534 719 820 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02533 1814 719 653 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02532 1814 716 1018 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02531 1018 716 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02530 718 722 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02529 730 893 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02528 655 728 729 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02527 1814 1173 655 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02526 830 729 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02525 1814 693 690 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02524 690 689 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02523 1814 711 689 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02522 1814 707 651 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02521 651 1173 650 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02520 650 706 709 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02519 708 709 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02518 1814 708 794 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02517 794 703 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02516 1814 878 703 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02515 759 707 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02514 648 759 693 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02513 1814 1708 648 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02512 1814 694 698 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02511 874 698 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02510 1814 701 698 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02509 698 695 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02508 1814 680 679 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02507 644 788 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02506 644 683 680 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02505 680 690 644 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02504 649 890 700 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02503 1814 759 649 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02502 701 700 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02501 1814 761 779 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02500 779 890 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02499 1814 685 779 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02498 779 1245 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02497 647 890 862 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02496 1814 1003 647 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02495 1814 681 645 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02494 645 682 646 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02493 646 862 684 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02492 683 684 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02491 640 995 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02490 660 671 640 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02489 662 672 660 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02488 666 672 642 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02487 642 662 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02486 641 671 666 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02485 672 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02484 1814 672 671 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02483 664 673 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02482 1814 664 641 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02481 1814 660 995 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02480 995 660 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02479 662 666 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02478 1814 670 643 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02477 673 679 643 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02476 643 675 673 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02475 1814 788 675 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02474 675 995 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02473 675 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02472 1814 623 624 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02471 626 624 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02470 1814 1245 624 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02469 624 833 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02468 1814 740 629 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02467 635 741 629 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02466 629 628 635 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02465 630 1245 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02464 631 638 630 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02463 632 639 631 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02462 634 639 633 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02461 633 632 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02460 636 638 634 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02459 639 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02458 1814 639 638 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02457 637 635 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02456 1814 637 636 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02455 1814 631 1245 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02454 1245 631 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02453 632 634 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02452 627 625 628 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02451 1814 626 627 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02450 625 908 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02449 1814 622 625 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02448 620 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02447 619 1325 621 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02446 1814 1244 619 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02445 621 618 620 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02444 617 621 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02443 761 1018 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02442 623 1239 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02441 1814 761 623 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02440 615 611 614 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02439 616 612 615 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02438 613 890 616 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02437 1814 618 613 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02436 1814 614 610 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02435 608 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02434 607 1201 609 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02433 1814 1244 607 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02432 609 612 608 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02431 606 609 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02430 707 601 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02429 1814 1086 707 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02428 1814 995 603 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02427 605 610 604 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02426 604 602 706 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02425 603 1003 605 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02424 1814 1003 597 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02423 600 610 599 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02422 599 602 598 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02421 597 596 600 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02420 694 1169 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02419 1814 598 694 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02418 589 1243 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02417 591 1115 590 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02416 1814 1244 591 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02415 590 588 589 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02414 587 590 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02413 1814 681 594 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02412 594 890 593 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02411 593 595 592 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02410 695 592 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02409 581 596 585 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02408 1814 995 581 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02407 681 585 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02406 1814 1708 583 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02405 583 601 584 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02404 584 595 586 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02403 582 586 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02402 577 1169 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02401 1814 577 579 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02400 579 578 601 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02399 580 1245 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02398 1814 761 580 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02397 1814 576 578 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02396 578 1239 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02395 1814 750 578 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02394 578 685 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02393 576 580 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02392 575 750 574 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02391 1814 1007 575 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02390 565 564 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02389 566 573 565 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02388 567 572 566 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02387 571 572 570 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02386 570 567 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02385 568 573 571 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02384 572 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02383 1814 572 573 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02382 569 606 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02381 1814 569 568 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02380 1814 566 564 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02379 564 566 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02378 567 571 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02377 685 1007 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02376 1814 553 472 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02375 472 560 473 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02374 473 557 555 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02373 554 555 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02372 1814 618 474 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02371 474 560 475 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02370 475 559 562 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02369 561 562 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02368 471 611 559 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02367 1814 612 471 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02366 470 549 550 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02365 1814 1708 470 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02364 551 550 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02363 549 546 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02362 1814 731 546 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02361 557 559 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02360 1814 612 461 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02359 463 602 462 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02358 462 521 523 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02357 461 878 463 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02356 1814 526 622 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02355 622 523 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02354 622 522 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02353 469 728 545 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02352 467 551 469 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02351 468 1007 467 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02350 1814 965 468 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02349 1814 545 560 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02348 833 1173 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02347 526 527 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02346 527 595 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02345 1814 588 527 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02344 527 711 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02343 1814 553 527 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02342 464 532 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02341 534 541 464 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02340 533 542 534 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02339 538 542 466 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02338 466 533 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02337 465 541 538 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02336 542 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02335 1814 542 541 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02334 536 617 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02333 1814 536 465 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02332 1814 534 532 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02331 532 534 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02330 533 538 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02329 1814 995 458 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02328 458 1173 459 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02327 459 878 516 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02326 514 516 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02325 508 512 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02324 512 819 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02323 1814 801 512 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02322 512 995 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02321 1814 1086 512 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02320 519 1086 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02319 1814 1169 519 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02318 518 833 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02317 1814 518 460 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02316 460 519 522 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02315 1814 506 502 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02314 502 1003 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02313 502 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02312 1814 500 501 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02311 456 506 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02310 456 582 500 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02309 500 498 456 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02308 455 1003 491 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02307 1814 682 455 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02306 498 491 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02305 1814 508 506 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02304 506 505 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02303 1814 1173 505 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02302 1814 670 457 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02301 503 501 457 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02300 457 502 503 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02299 449 580 487 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02298 450 728 449 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02297 451 488 450 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02296 1814 574 451 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02295 1814 487 484 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02294 476 478 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02293 1814 532 478 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02292 452 728 490 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02291 453 489 452 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02290 454 965 453 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02289 1814 488 454 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02288 1814 490 682 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02287 479 477 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02286 1814 848 477 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02285 1814 484 482 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02284 482 481 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02283 1814 596 481 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02282 1814 670 437 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02281 438 440 437 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02280 437 439 438 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02279 1814 448 446 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02278 447 445 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02277 447 561 448 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02276 448 444 447 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02275 1814 445 439 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02274 439 612 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02273 439 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02272 428 612 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02271 430 436 428 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02270 431 434 430 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02269 433 434 432 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02268 432 431 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02267 429 436 433 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02266 434 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02265 1814 434 436 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02264 435 438 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02263 1814 435 429 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02262 1814 430 612 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02261 612 430 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02260 431 433 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02259 1814 443 440 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02258 442 445 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02257 442 554 443 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02256 443 441 442 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02255 1814 521 444 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02254 444 618 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02253 444 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02252 553 618 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02251 1814 965 426 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02250 426 1007 425 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02249 425 731 427 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02248 424 427 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02247 423 915 422 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02246 1814 622 423 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02245 421 422 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02244 420 1086 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02243 1814 595 420 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02242 1814 801 414 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02241 414 711 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02240 414 1015 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02239 878 801 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02238 1814 1173 416 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02237 416 420 418 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02236 418 417 419 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02235 415 419 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02234 1814 801 417 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02233 417 711 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02232 417 1015 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02231 596 1086 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02230 404 415 403 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02229 1814 400 404 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02228 402 403 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02227 405 1003 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02226 406 412 405 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02225 407 413 406 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02224 409 413 408 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02223 408 407 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02222 410 412 409 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02221 413 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02220 1814 413 412 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02219 411 503 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02218 1814 411 410 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02217 1814 406 1003 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02216 1003 406 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02215 407 409 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02214 398 1086 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02213 1814 1173 398 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02212 375 1086 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02211 374 382 375 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02210 373 381 374 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02209 377 381 379 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02208 379 373 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02207 378 382 377 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02206 381 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02205 1814 381 382 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02204 376 396 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02203 1814 376 378 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02202 1814 374 1086 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02201 1086 374 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02200 373 377 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02199 1814 391 397 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02198 396 395 397 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02197 397 399 396 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02196 1814 398 401 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02195 399 401 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02194 1814 402 401 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02193 401 908 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02192 380 965 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02191 1814 384 380 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02190 386 576 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02189 1814 1007 386 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02188 385 386 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02187 1814 385 383 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02186 383 1708 384 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02185 1814 393 395 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02184 394 1173 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02183 394 482 393 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02182 393 392 394 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02181 387 386 390 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02180 388 728 387 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02179 389 1086 388 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02178 1814 488 389 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02177 1814 390 392 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02176 1814 670 292 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02175 363 446 292 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02174 292 361 363 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02173 243 618 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02172 365 297 243 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02171 368 298 365 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02170 367 298 295 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02169 295 368 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02168 294 297 367 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02167 298 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02166 1814 298 297 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02165 296 363 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02164 1814 296 294 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02163 1814 365 618 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02162 618 365 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02161 368 367 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02160 291 915 356 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02159 1814 333 291 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02158 445 356 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02157 1814 445 361 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02156 361 618 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02155 361 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02154 350 612 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02153 346 345 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02152 1814 424 345 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02151 1814 351 341 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02150 341 1086 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02149 1814 337 341 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02148 341 595 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02147 1814 612 290 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02146 290 618 289 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02145 289 611 349 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02144 351 349 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02143 1814 893 347 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02142 347 553 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02141 347 350 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02140 286 488 343 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02139 287 346 286 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02138 288 351 287 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02137 1814 415 288 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02136 1814 343 344 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02135 1814 965 278 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02134 278 279 280 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02133 280 347 328 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02132 400 328 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02131 282 1086 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02130 1814 595 282 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02129 595 1003 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02128 279 588 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02127 1814 685 279 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02126 283 414 331 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02125 284 488 283 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02124 285 1173 284 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02123 1814 282 285 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02122 1814 331 333 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02121 1814 322 391 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02120 276 1708 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02119 276 915 322 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02118 322 596 276 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02117 266 685 267 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02116 1814 1708 266 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02115 1814 400 274 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02114 274 415 275 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02113 275 488 325 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02112 326 325 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02111 189 300 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02110 301 258 189 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02109 303 259 301 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02108 302 259 255 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02107 255 303 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02106 254 258 302 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02105 259 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02104 1814 259 258 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02103 256 587 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02102 1814 256 254 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02101 1814 301 300 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02100 300 301 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02099 303 302 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02098 270 915 317 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02097 271 272 270 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02096 269 596 271 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02095 1814 1173 269 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02094 1814 317 319 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02093 272 268 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02092 1814 319 312 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02091 312 965 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02090 312 1758 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02089 1814 308 309 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02088 260 319 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02087 260 380 308 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02086 308 315 260 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02085 265 576 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02084 1814 1758 265 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02083 1814 265 263 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02082 263 965 262 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02081 262 685 313 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02080 315 313 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02079 1814 234 233 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02078 235 1708 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02077 235 915 234 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02076 234 611 235 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02075 611 588 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02074 1814 1708 241 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02073 241 350 239 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02072 239 238 240 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02071 441 240 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02070 238 237 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02069 1814 588 237 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02068 237 236 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02067 242 819 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02066 247 252 242 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02065 244 250 247 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02064 246 250 245 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02063 245 244 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02062 249 252 246 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02061 250 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02060 1814 250 252 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02059 251 248 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02058 1814 251 249 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02057 1814 247 819 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02056 819 247 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02055 244 246 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02054 521 231 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02053 1814 230 231 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02052 232 230 236 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02051 1814 553 232 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02050 230 229 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02049 228 424 229 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02048 1814 728 228 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02047 337 227 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02046 1814 229 227 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02045 1814 1015 226 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02044 225 488 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02043 226 341 225 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02042 670 224 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02041 1814 1003 220 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02040 221 1015 222 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02039 222 521 223 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02038 220 596 221 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02037 1814 217 216 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02036 218 514 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02035 218 226 217 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02034 217 219 218 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02033 219 1169 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02032 1814 223 219 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02031 213 214 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02030 1814 1007 214 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02029 214 215 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02028 208 576 215 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02027 1814 1708 208 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02026 202 204 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02025 207 203 205 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02024 207 272 1814 1814 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02023 1814 267 207 1814 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02022 205 213 204 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02021 204 268 207 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02020 268 206 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02019 1814 1169 206 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02018 206 1239 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02017 1814 965 209 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02016 211 728 210 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02015 210 215 212 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02014 209 596 211 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02013 203 489 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02012 200 1007 201 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02011 1814 265 200 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02010 489 201 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02009 186 187 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02008 1814 300 187 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02007 1814 670 199 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02006 198 309 199 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02005 199 312 198 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02004 188 965 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02003 193 196 188 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02002 190 197 193 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02001 192 197 191 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02000 191 190 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01999 195 196 192 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01998 197 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01997 1814 197 196 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01996 194 198 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01995 1814 194 195 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01994 1814 193 965 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01993 965 193 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01992 190 192 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01991 160 155 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01990 1814 588 162 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01989 158 160 156 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01988 156 588 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01987 156 162 158 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01986 1814 155 156 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01985 161 166 248 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01984 1814 1708 161 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01983 155 154 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01982 1814 236 154 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01981 138 137 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01980 1814 1239 137 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01979 137 908 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01978 1814 163 164 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01977 164 165 166 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01976 164 819 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01975 166 184 164 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01974 1814 819 165 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01973 163 184 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01972 1814 143 141 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01971 64 1708 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01970 64 915 143 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01969 143 728 64 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01968 602 1015 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01967 1814 141 140 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01966 146 344 140 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01965 140 138 146 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01964 1814 1708 133 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01963 134 421 133 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01962 133 132 134 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01961 66 1239 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01960 145 153 66 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01959 147 152 145 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01958 150 152 69 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01957 69 147 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01956 68 153 150 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01955 152 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01954 1814 152 153 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01953 149 146 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01952 1814 149 68 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01951 1814 145 1239 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01950 1239 145 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01949 147 150 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01948 47 1015 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01947 114 120 47 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01946 115 121 114 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01945 118 121 50 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01944 50 115 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01943 49 120 118 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01942 121 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01941 1814 121 120 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01940 119 127 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01939 1814 119 49 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01938 1814 114 1015 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01937 1015 114 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01936 115 118 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01935 1814 128 126 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01934 127 216 126 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01933 126 125 127 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01932 103 915 105 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01931 1814 1173 103 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01930 1814 122 123 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01929 125 1015 123 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01928 123 514 125 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01927 1814 131 128 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01926 53 1708 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01925 53 915 131 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01924 131 602 53 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01923 112 1169 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01922 1814 212 112 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01921 99 267 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01920 1814 99 100 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01919 100 105 102 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01918 1814 98 96 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01917 98 224 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01916 1814 101 36 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01915 36 102 98 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01914 1814 202 104 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01913 101 104 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01912 1814 105 104 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01911 104 112 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01910 1814 109 108 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01909 44 1708 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01908 44 915 109 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01907 109 488 44 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01906 728 1239 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01905 23 1007 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01904 86 91 23 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01903 85 92 86 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01902 88 92 27 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01901 27 85 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01900 26 91 88 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01899 92 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01898 1814 92 91 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01897 87 96 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01896 1814 87 26 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01895 1814 86 1007 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01894 1007 86 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01893 85 88 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01892 95 94 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01891 1814 1239 94 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01890 94 576 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01889 1814 65 67 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01888 70 588 67 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01887 67 333 70 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01886 74 588 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01885 78 83 74 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01884 75 81 78 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01883 77 81 76 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01882 76 75 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01881 80 83 77 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01880 81 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01879 1814 81 83 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01878 82 79 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01877 1814 82 80 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01876 1814 78 588 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01875 588 78 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01874 75 77 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01873 1814 233 71 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01872 79 73 71 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01871 71 70 79 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01870 65 908 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01869 1814 158 73 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01868 73 72 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01867 1814 333 72 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01866 132 54 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01865 55 54 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01864 56 62 55 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01863 57 63 56 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01862 59 63 60 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01861 60 57 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01860 58 62 59 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01859 63 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01858 1814 63 62 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01857 61 134 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01856 1814 61 58 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01855 1814 56 54 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01854 54 56 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01853 57 59 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01852 52 819 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01851 1814 52 51 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01850 51 54 908 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01849 224 54 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01848 1814 819 224 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01847 488 1169 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01846 122 908 1814 1814 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01845 1814 326 46 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01844 45 46 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01843 1814 908 46 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01842 46 48 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01841 1814 108 43 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01840 42 45 43 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01839 43 41 42 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01838 25 1169 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01837 24 34 25 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01836 28 33 24 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01835 30 33 31 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01834 31 28 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01833 29 34 30 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01832 33 1810 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01831 1814 33 34 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01830 32 42 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01829 1814 32 29 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01828 1814 24 1169 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01827 1169 24 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01826 28 30 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01825 48 1169 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01824 1814 1173 48 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01823 35 1169 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01822 1814 95 37 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01821 39 35 38 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01820 38 95 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01819 38 37 39 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01818 1814 1169 38 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01817 1814 39 41 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01816 41 40 1814 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01815 1814 1173 40 1814 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01814 22 21 1814 1814 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01813 1814 564 21 1814 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01812 1727 1793 1706 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01811 1706 1792 1795 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01810 1795 1791 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01809 1727 1801 1802 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01808 1727 1798 1809 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01807 1727 1796 1713 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01806 1713 1795 1727 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01805 1798 1802 1712 1727 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01804 1712 1808 1727 1727 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01803 1713 1797 1798 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01802 1788 1808 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01801 1727 1786 1787 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01800 1703 1787 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01799 1797 1788 1703 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01798 1702 1786 1797 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01797 1727 1808 1702 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01796 1718 1815 1804 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01795 1727 1808 1718 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01794 1804 1813 1805 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01793 1727 1805 1723 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01792 1723 1813 1807 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01791 1807 1815 1725 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01790 1813 1815 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01789 1727 1810 1815 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01788 1725 1812 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01787 1727 1809 1812 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01786 1808 1804 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01785 1727 1804 1808 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01784 1805 1807 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01783 1784 1780 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01782 1727 1778 1784 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01781 1775 1771 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01780 1775 1778 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01779 1727 1772 1775 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01778 1727 1775 1790 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01777 1727 1784 1699 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01776 1699 1785 1698 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01775 1698 1783 1793 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01774 1777 1786 1691 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01773 1727 1777 1780 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01772 1691 1776 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01771 1782 1780 1694 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01770 1727 1782 1781 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01769 1694 1792 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01768 1727 1769 1685 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01767 1685 1783 1770 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01766 1759 1761 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01765 1727 1765 1761 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01764 1671 1764 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01763 1761 1771 1671 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01762 1727 1768 1765 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01761 1679 1770 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01760 1680 1785 1679 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01759 1768 1767 1680 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01758 1676 1772 1764 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01757 1764 1766 1676 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01756 1676 1762 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01755 1727 1767 1766 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01754 1755 1769 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01753 1727 1752 1754 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01752 1662 1754 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01751 1757 1755 1662 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01750 1663 1752 1757 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01749 1727 1769 1663 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01748 1727 1758 1668 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01747 1668 1772 1669 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01746 1669 1757 1762 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01745 1653 1753 1746 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01744 1727 1752 1653 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01743 1746 1748 1747 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01742 1727 1747 1652 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01741 1652 1748 1751 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01740 1751 1753 1656 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01739 1748 1753 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01738 1727 1810 1753 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01737 1656 1749 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01736 1727 1759 1749 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01735 1752 1746 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01734 1727 1746 1752 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01733 1747 1751 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01732 1727 1743 1742 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01731 1647 1785 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01730 1648 1772 1647 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01729 1743 1758 1648 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01728 1632 1737 1730 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01727 1727 1772 1632 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01726 1730 1738 1731 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01725 1727 1731 1637 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01724 1637 1738 1735 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01723 1735 1737 1638 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01722 1738 1737 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01721 1727 1810 1737 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01720 1638 1733 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01719 1727 1736 1733 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01718 1772 1730 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01717 1727 1730 1772 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01716 1731 1735 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01715 1736 1741 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01714 1727 1742 1741 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01713 1645 1739 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01712 1741 1771 1645 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01711 1714 1790 1801 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01710 1801 1710 1714 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01709 1714 1758 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01708 1727 1722 1717 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01707 1717 1715 1796 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01706 1796 1716 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01705 1704 1790 1705 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01704 1727 1704 1707 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01703 1705 1792 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01702 1722 1721 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01701 1727 1726 1721 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01700 1720 1719 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01699 1721 1776 1720 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01698 1711 1707 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01697 1711 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01696 1727 1709 1711 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01695 1727 1711 1716 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01694 1727 1808 1792 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01693 1697 1695 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01692 1697 1772 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01691 1727 1701 1697 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01690 1727 1697 1696 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01689 1726 1724 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01688 1724 1772 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01687 1727 1771 1724 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01686 1693 1778 1692 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01685 1727 1693 1695 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01684 1692 1776 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01683 1727 1758 1700 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01682 1700 1785 1701 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01681 1727 1655 1657 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01680 1655 1654 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01679 1727 1771 1785 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01678 1727 1772 1783 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01677 1660 1657 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01676 1727 1786 1658 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01675 1661 1658 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01674 1664 1660 1661 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01673 1659 1786 1664 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01672 1727 1657 1659 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01671 1767 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01670 1727 1677 1767 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01669 1678 1690 1686 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01668 1727 1786 1678 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01667 1686 1689 1681 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01666 1727 1681 1682 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01665 1682 1689 1684 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01664 1684 1690 1683 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01663 1689 1690 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01662 1727 1810 1690 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01661 1683 1688 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01660 1727 1687 1688 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01659 1786 1686 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01658 1727 1686 1786 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01657 1681 1684 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01656 1674 1672 1675 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01655 1727 1674 1673 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01654 1675 1758 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01653 1666 1664 1665 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01652 1727 1673 1666 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01651 1667 1670 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01650 1665 1786 1667 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01649 1727 1665 1687 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01648 1670 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01647 1727 1672 1670 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01646 1727 1646 1643 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01645 1643 1772 1644 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01644 1727 1772 1649 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01643 1644 1649 1642 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01642 1642 1641 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01641 1739 1644 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01640 1646 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01639 1727 1769 1646 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01638 1727 1651 1769 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01637 1651 1650 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01636 1631 1639 1630 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01635 1727 1650 1631 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01634 1630 1640 1629 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01633 1727 1629 1634 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01632 1634 1640 1635 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01631 1635 1639 1636 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01630 1640 1639 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01629 1727 1810 1639 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01628 1636 1633 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01627 1727 1646 1633 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01626 1650 1630 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01625 1727 1630 1650 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01624 1629 1635 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01623 1719 1603 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01622 1603 1602 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01621 1727 1601 1603 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01620 1596 1592 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01619 1592 1696 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01618 1727 1709 1592 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01617 1606 1808 1551 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01616 1727 1606 1715 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01615 1551 1605 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01614 1727 1776 1540 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01613 1540 1600 1598 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01612 1598 1596 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01611 1599 1602 1541 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01610 1727 1599 1600 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01609 1541 1715 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01608 1727 1710 1585 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01607 1727 1586 1529 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01606 1529 1585 1587 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01605 1594 1595 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01604 1595 1808 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01603 1727 1776 1595 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01602 1727 1696 1590 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01601 1590 1587 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01600 1590 1781 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01599 1778 1583 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01598 1583 1601 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01597 1727 1582 1583 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01596 1727 1579 1509 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01595 1509 1710 1578 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01594 1727 1580 1579 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01593 1511 1783 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01592 1512 1785 1511 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01591 1580 1581 1512 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01590 1577 1579 1507 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01589 1727 1577 1672 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01588 1507 1585 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01587 1727 1581 1601 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01586 1727 1654 1582 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01585 1727 1565 1564 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01584 1490 1567 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01583 1494 1785 1490 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01582 1565 1641 1494 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01581 1727 1576 1677 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01580 1576 1575 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01579 1654 1575 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01578 1727 1574 1654 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01577 1727 1570 1654 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01576 1654 1569 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01575 1727 1650 1570 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01574 1567 1568 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01573 1568 1772 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01572 1727 1677 1568 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01571 1727 1752 1575 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01570 1562 1561 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01569 1727 1564 1561 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01568 1488 1771 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01567 1561 1646 1488 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01566 1478 1558 1552 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01565 1727 1771 1478 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01564 1552 1560 1554 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01563 1727 1554 1483 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01562 1483 1560 1556 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01561 1556 1558 1482 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01560 1560 1558 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01559 1727 1810 1558 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01558 1482 1559 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01557 1727 1562 1559 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01556 1771 1552 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01555 1727 1552 1771 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01554 1554 1556 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01553 1537 1792 1538 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01552 1538 1535 1537 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01551 1537 1594 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01550 1727 1543 1534 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01549 1534 1531 1535 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01548 1535 1532 1533 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01547 1533 1786 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01546 1727 1786 1531 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01545 1532 1543 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01544 1727 1801 1468 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01543 1727 1539 1550 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01542 1727 1590 1467 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01541 1467 1598 1727 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01540 1539 1468 1466 1727 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01539 1466 1543 1727 1727 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01538 1467 1538 1539 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01537 1470 1548 1542 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01536 1727 1543 1470 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01535 1542 1545 1547 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01534 1727 1547 1546 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01533 1546 1545 1544 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01532 1544 1548 1473 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01531 1545 1548 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01530 1727 1810 1548 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01529 1473 1549 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01528 1727 1550 1549 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01527 1543 1542 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01526 1727 1542 1543 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01525 1547 1544 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01524 1727 1776 1522 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01523 1522 1792 1521 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01522 1521 1585 1520 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01521 1727 1783 1525 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01520 1525 1785 1527 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01519 1527 1523 1526 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01518 1526 1524 1528 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01517 1523 1530 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01516 1727 1710 1523 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01515 1727 1594 1463 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01514 1463 1536 1530 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01513 1727 1808 1459 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01512 1459 1776 1524 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01511 1727 1502 1505 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01510 1505 1585 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01509 1519 1501 1505 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01508 1505 1506 1519 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01507 1506 1503 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01506 1503 1508 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01505 1727 1504 1503 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01504 1727 1581 1497 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01503 1501 1497 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01502 1727 1569 1501 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01501 1453 1581 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01500 1727 1508 1453 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01499 1727 1771 1453 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01498 1453 1585 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01497 1455 1518 1510 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01496 1727 1710 1455 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01495 1510 1513 1517 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01494 1727 1517 1516 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01493 1516 1513 1515 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01492 1515 1518 1458 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01491 1513 1518 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01490 1727 1810 1518 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01489 1458 1514 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01488 1727 1519 1514 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01487 1710 1510 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01486 1727 1510 1710 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01485 1517 1515 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01484 1508 1499 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01483 1499 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01482 1727 1500 1499 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01481 1641 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01480 1727 1570 1641 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01479 1727 1498 1500 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01478 1442 1677 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01477 1727 1570 1442 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01476 1727 1677 1498 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01475 1498 1574 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01474 1498 1570 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01473 1439 1495 1486 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01472 1727 1489 1439 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01471 1436 1485 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01470 1486 1578 1436 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01469 1727 1486 1487 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01468 1489 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01467 1727 1578 1489 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01466 1492 1498 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01465 1727 1569 1491 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01464 1493 1491 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01463 1495 1492 1493 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01462 1496 1569 1495 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01461 1727 1498 1496 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01460 1431 1484 1475 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01459 1727 1569 1431 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01458 1475 1479 1477 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01457 1727 1477 1481 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01456 1481 1479 1476 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01455 1476 1484 1434 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01454 1479 1484 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01453 1727 1810 1484 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01452 1434 1480 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01451 1727 1487 1480 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01450 1569 1475 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01449 1727 1475 1569 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01448 1477 1476 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01447 1415 1409 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01446 1727 1414 1415 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01445 1412 1410 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01444 1412 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01443 1727 1710 1412 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01442 1727 1412 1791 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01441 1727 1543 1776 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01440 1414 1419 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01439 1419 1601 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01438 1727 1417 1419 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01437 1406 1408 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01436 1408 1709 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01435 1727 1414 1408 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01434 1340 1428 1421 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01433 1727 1586 1340 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01432 1421 1429 1422 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01431 1727 1422 1342 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01430 1342 1429 1424 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01429 1424 1428 1343 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01428 1429 1428 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01427 1727 1810 1428 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01426 1343 1426 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01425 1727 1425 1426 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01424 1586 1421 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01423 1727 1421 1586 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01422 1422 1424 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01421 1727 1776 1336 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01420 1336 1415 1335 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01419 1335 1785 1332 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01418 1332 1783 1405 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01417 1403 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01416 1727 1410 1403 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01415 1400 1771 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01414 1727 1792 1400 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01413 1727 1406 1400 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01412 1400 1776 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01411 1330 1403 1402 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01410 1727 1528 1330 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01409 1331 1400 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01408 1402 1783 1331 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01407 1727 1402 1425 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01406 1379 1504 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01405 1318 1485 1382 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01404 1727 1379 1318 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01403 1727 1502 1321 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01402 1321 1601 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01401 1384 1601 1321 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01400 1321 1382 1384 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01399 1324 1396 1388 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01398 1727 1581 1324 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01397 1388 1395 1387 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01396 1727 1387 1327 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01395 1327 1395 1394 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01394 1394 1396 1328 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01393 1395 1396 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01392 1727 1810 1396 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01391 1328 1391 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01390 1727 1390 1391 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01389 1581 1388 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01388 1727 1388 1581 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01387 1387 1394 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01386 1390 1386 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01385 1727 1384 1386 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01384 1323 1453 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01383 1386 1783 1323 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01382 1727 1785 1320 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01381 1320 1783 1380 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01380 1727 1376 1312 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01379 1312 1758 1375 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01378 1316 1500 1502 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01377 1502 1380 1316 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01376 1316 1758 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01375 1299 1360 1351 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01374 1727 1349 1299 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01373 1351 1357 1350 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01372 1727 1350 1301 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01371 1301 1357 1356 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01370 1356 1360 1302 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01369 1357 1360 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01368 1727 1810 1360 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01367 1302 1354 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01366 1727 1353 1354 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01365 1349 1351 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01364 1727 1351 1349 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01363 1350 1356 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01362 1374 1574 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01361 1374 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01360 1727 1376 1374 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01359 1727 1374 1370 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01358 1727 1380 1376 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01357 1727 1347 1474 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01356 1347 1359 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01355 1727 1348 1728 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01354 1348 1349 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01353 1304 1371 1363 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01352 1727 1359 1304 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01351 1363 1369 1361 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01350 1727 1361 1305 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01349 1305 1369 1368 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01348 1368 1371 1309 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01347 1369 1371 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01346 1727 1810 1371 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01345 1309 1366 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01344 1727 1365 1366 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01343 1359 1363 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01342 1727 1363 1359 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01341 1361 1368 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01340 1727 1346 1345 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01339 1346 1344 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01338 1377 1758 1315 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01337 1727 1377 1485 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01336 1315 1569 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01335 1334 1333 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01334 1282 1334 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01333 1727 1334 1282 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01332 1727 1334 1282 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01331 1282 1334 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01330 1536 1601 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01329 1727 1282 1536 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01328 1727 1326 1605 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01327 1339 1605 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01326 1727 1601 1339 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01325 1727 1325 1339 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01324 1339 1417 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01323 1293 1339 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01322 1409 1341 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01321 1341 1326 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01320 1727 1808 1341 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01319 1727 1409 1289 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01318 1289 1536 1288 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01317 1276 1808 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01316 1727 1771 1276 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01315 1285 1337 1286 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01314 1286 1338 1285 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01313 1285 1405 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01312 1727 1329 1338 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01311 1278 1281 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01310 1277 1276 1278 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01309 1329 1783 1277 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01308 1727 1758 1287 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01307 1287 1326 1337 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01306 1727 1601 1281 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01305 1281 1282 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01304 1281 1543 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01303 1319 1267 1266 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01302 1727 1319 1265 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01301 1266 1758 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01300 1727 1708 1758 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01299 1322 1271 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01298 1727 1520 1322 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01297 1727 1772 1322 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01296 1322 1771 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01295 1267 1322 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01294 1727 1586 1273 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01293 1273 1325 1274 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01292 1274 1326 1272 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01291 1272 1581 1271 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01290 1317 1771 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01289 1317 1710 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01288 1727 1772 1317 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01287 1727 1317 1504 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01286 1255 1264 1311 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01285 1727 1308 1255 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01284 1311 1259 1313 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01283 1727 1313 1256 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01282 1256 1259 1314 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01281 1314 1264 1261 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01280 1259 1264 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01279 1727 1810 1264 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01278 1261 1260 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01277 1727 1257 1260 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01276 1308 1311 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01275 1727 1311 1308 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01274 1313 1314 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01273 1727 1442 1250 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01272 1250 1306 1310 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01271 1310 1307 1251 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01270 1251 1308 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01269 1727 1308 1306 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01268 1307 1442 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01267 1242 1769 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01266 1727 1244 1242 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01265 1242 1243 1300 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01264 1300 1239 1242 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01263 1727 1300 1353 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01262 1253 1375 1257 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01261 1257 1310 1253 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01260 1253 1370 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01259 1248 1245 1303 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01258 1727 1244 1248 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01257 1247 1243 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01256 1303 1752 1247 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01255 1727 1303 1241 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01254 1727 1295 1228 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01253 1295 1229 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01252 1230 1238 1296 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01251 1727 1344 1230 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01250 1296 1235 1297 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01249 1727 1297 1232 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01248 1232 1235 1298 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01247 1298 1238 1236 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01246 1235 1238 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01245 1727 1810 1238 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01244 1236 1234 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01243 1727 1241 1234 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01242 1344 1296 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01241 1727 1296 1344 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01240 1297 1298 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01239 1150 1219 1213 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01238 1727 1326 1150 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01237 1213 1220 1214 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01236 1727 1214 1151 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01235 1151 1220 1216 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01234 1216 1219 1152 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01233 1220 1219 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01232 1727 1810 1219 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01231 1152 1218 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01230 1727 1221 1218 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01229 1326 1213 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01228 1727 1213 1326 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01227 1214 1216 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01226 1727 1225 1226 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01225 1727 1227 1224 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01224 1154 1226 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01223 1155 1326 1154 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01222 1227 1758 1155 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01221 1417 1211 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01220 1211 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01219 1727 1333 1211 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01218 1221 1222 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01217 1727 1224 1222 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01216 1153 1286 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01215 1222 1225 1153 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01214 1207 1204 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01213 1727 1582 1207 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01212 1727 1206 1208 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01211 1727 1207 1333 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01210 1203 1201 1147 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01209 1727 1203 1202 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01208 1147 1204 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01207 1727 1786 1204 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01206 1727 1209 1602 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01205 1149 1208 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01204 1148 1786 1149 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01203 1209 1325 1148 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01202 1144 1198 1192 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01201 1727 1190 1144 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01200 1192 1199 1194 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01199 1727 1194 1145 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01198 1145 1199 1196 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01197 1196 1198 1146 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01196 1199 1198 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01195 1727 1810 1198 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01194 1146 1200 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01193 1727 1193 1200 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01192 1190 1192 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01191 1727 1192 1190 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01190 1194 1196 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01189 1186 1185 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01188 1727 1201 1184 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01187 1142 1184 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01186 1188 1186 1142 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01185 1141 1201 1188 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01184 1727 1185 1141 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01183 1189 1188 1143 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01182 1727 1189 1187 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01181 1143 1786 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01180 1185 1569 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01179 1727 1178 1185 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01178 1727 1574 1185 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01177 1185 1177 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01176 1727 1308 1574 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01175 1140 1173 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01174 1727 1243 1140 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01173 1140 1244 1176 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01172 1176 1772 1140 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01171 1727 1176 1365 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01170 1139 1308 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01169 1727 1244 1139 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01168 1139 1243 1171 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01167 1171 1169 1139 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01166 1727 1171 1167 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01165 1727 1442 1178 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01164 1137 1168 1162 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01163 1727 1229 1137 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01162 1162 1163 1160 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01161 1727 1160 1136 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01160 1136 1163 1165 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01159 1165 1168 1138 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01158 1163 1168 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01157 1727 1810 1168 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01156 1138 1164 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01155 1727 1167 1164 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01154 1229 1162 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01153 1727 1162 1229 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01152 1160 1165 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01151 1727 1156 1157 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01150 1156 1190 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01149 1727 1808 1126 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01148 1126 1206 1127 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01147 1128 1288 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01146 1727 1710 1128 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01145 1727 1771 1133 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01144 1133 1543 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01143 1133 1772 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01142 1727 1134 1130 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01141 1130 1128 1132 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01140 1132 1133 1131 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01139 1131 1127 1129 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01138 1727 1326 1135 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01137 1135 1808 1134 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01136 1727 1586 1410 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01135 1090 1201 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01134 1089 1177 1206 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01133 1727 1090 1089 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01132 1727 1113 1114 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01131 1113 1207 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01130 1112 1114 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01129 1727 1115 1108 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01128 1109 1108 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01127 1110 1112 1109 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01126 1111 1115 1110 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01125 1727 1114 1111 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01124 1727 1115 1177 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01123 1116 1125 1118 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01122 1727 1115 1116 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01121 1118 1124 1117 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01120 1727 1117 1120 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01119 1120 1124 1119 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01118 1119 1125 1121 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01117 1124 1125 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01116 1727 1810 1125 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01115 1121 1123 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01114 1727 1122 1123 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01113 1115 1118 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01112 1727 1118 1115 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01111 1117 1119 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01110 1104 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01109 1727 1267 1104 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01108 1727 1103 1100 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01107 1727 1187 1101 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01106 1101 1202 1727 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01105 1103 1265 1102 1727 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01104 1102 1201 1727 1727 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01103 1101 1104 1103 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01102 1091 1098 1092 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01101 1727 1201 1091 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01100 1092 1097 1093 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01099 1727 1093 1094 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01098 1094 1097 1095 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01097 1095 1098 1096 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01096 1097 1098 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01095 1727 1810 1098 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01094 1096 1099 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01093 1727 1100 1099 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01092 1201 1092 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01091 1727 1092 1201 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01090 1093 1095 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01089 1107 1110 1106 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01088 1727 1104 1107 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01087 1105 1265 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01086 1106 1115 1105 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01085 1727 1106 1122 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01084 1088 1581 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01083 1727 1244 1088 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01082 1088 1243 1087 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01081 1087 1086 1088 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01080 1727 1087 1085 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01079 1074 1084 1076 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01078 1727 1075 1074 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01077 1076 1083 1078 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01076 1727 1078 1081 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01075 1081 1083 1080 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01074 1080 1084 1082 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01073 1083 1084 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01072 1727 1810 1084 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01071 1082 1079 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01070 1727 1077 1079 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01069 1075 1076 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01068 1727 1076 1075 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01067 1078 1080 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01066 1065 1072 1066 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01065 1727 1064 1065 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01064 1066 1071 1067 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01063 1727 1067 1068 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01062 1068 1071 1070 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01061 1070 1072 1069 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01060 1071 1072 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01059 1727 1810 1072 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01058 1069 1073 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01057 1727 1085 1073 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01056 1064 1066 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01055 1727 1066 1064 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01054 1067 1070 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01053 1727 1062 1607 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01052 1062 1075 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01051 1727 1063 1061 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01050 1063 1064 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01049 1225 1710 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01048 1727 1410 1225 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01047 1043 1050 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01046 1727 1709 1043 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01045 1727 1326 947 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01044 947 1050 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01043 1052 1057 947 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01042 947 1293 1052 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01041 1042 1049 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01040 1727 1326 944 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01039 944 1043 1049 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01038 946 1047 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01037 1727 1044 945 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01036 1049 1052 946 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01035 945 1129 1049 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01034 1058 1772 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01033 1727 1771 1058 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01032 1727 1808 1058 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01031 1058 1543 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01030 1057 1058 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01029 1047 1710 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01028 1727 1410 1047 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01027 1709 1036 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01026 1036 1586 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01025 1727 1710 1036 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01024 941 1031 1024 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01023 1727 1173 941 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01022 1024 1033 1026 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01021 1727 1026 942 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01020 942 1033 1029 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01019 1029 1031 943 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01018 1033 1031 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01017 1727 1810 1031 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01016 943 1032 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01015 1727 1027 1032 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01014 1173 1024 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01013 1727 1024 1173 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01012 1026 1029 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01011 1727 1244 1243 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01010 940 1018 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01009 1727 1243 940 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01008 940 1244 1019 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01007 1019 1771 940 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01006 1727 1019 1077 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01005 936 995 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01004 1727 1243 936 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01003 936 1244 997 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01002 997 1808 936 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01001 1727 997 993 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01000 938 1710 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00999 1727 1244 938 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00998 938 1243 1010 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00997 1010 1007 938 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00996 1727 1010 1193 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00995 937 1003 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00994 1727 1243 937 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00993 937 1244 1004 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00992 1004 1543 937 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00991 1727 1004 1001 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00990 939 1326 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00989 1727 1244 939 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00988 939 1243 1016 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00987 1016 1015 939 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00986 1727 1016 1012 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00985 930 981 972 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00984 1727 969 930 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00983 972 978 971 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00982 1727 971 932 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00981 932 978 977 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00980 977 981 931 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00979 978 981 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00978 1727 1810 981 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00977 931 975 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00976 1727 993 975 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00975 969 972 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00974 1727 972 969 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00973 971 977 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00972 929 1569 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00971 1727 1244 929 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00970 929 1243 966 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00969 966 965 929 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00968 1727 966 962 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00967 934 992 985 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00966 1727 980 934 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00965 985 988 986 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00964 1727 986 933 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00963 933 988 991 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00962 991 992 935 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00961 988 992 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00960 1727 1810 992 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00959 935 989 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00958 1727 1012 989 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00957 980 985 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00956 1727 985 980 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00955 986 991 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00954 926 963 955 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00953 1727 950 926 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00952 955 959 952 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00951 1727 952 927 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00950 927 959 954 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00949 954 963 928 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00948 959 963 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00947 1727 1810 963 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00946 928 957 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00945 1727 962 957 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00944 950 955 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00943 1727 955 950 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00942 952 954 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00941 1727 948 949 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00940 948 950 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00939 917 925 920 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00938 1727 1325 917 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00937 920 924 921 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00936 1727 921 918 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00935 918 924 919 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00934 919 925 922 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00933 924 925 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00932 1727 1810 925 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00931 922 923 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00930 1727 1042 923 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00929 1325 920 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00928 1727 920 1325 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00927 921 919 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00926 914 1018 913 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00925 1727 914 912 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00924 913 1239 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00923 1727 1325 916 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00922 1044 916 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00921 1727 1708 1044 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00920 1727 1044 1050 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00919 1727 905 909 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00918 906 915 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00917 904 1173 906 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00916 905 1758 904 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00915 1727 908 880 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00914 896 903 895 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00913 1727 893 896 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00912 895 902 897 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00911 1727 897 894 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00910 894 902 900 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00909 900 903 901 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00908 902 903 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00907 1727 1810 903 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00906 901 899 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00905 1727 898 899 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00904 893 895 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00903 1727 895 893 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00902 897 900 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00901 1027 911 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00900 1727 909 911 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00899 910 907 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00898 911 908 910 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00897 892 1586 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00896 1727 1244 892 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00895 892 1243 891 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00894 891 893 892 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00893 1727 891 889 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00892 1727 893 882 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00891 882 881 884 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00890 884 880 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00889 881 879 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00888 879 1173 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00887 1727 878 879 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00886 1727 883 886 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00885 886 884 898 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00884 898 887 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00883 865 873 866 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00882 1727 864 865 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00881 866 872 867 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00880 1727 867 869 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00879 869 872 870 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00878 870 873 871 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00877 872 873 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00876 1727 1810 873 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00875 871 868 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00874 1727 1001 868 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00873 864 866 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00872 1727 866 864 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00871 867 870 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00870 887 885 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00869 1727 1708 885 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00868 888 915 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00867 885 890 888 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00866 883 877 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00865 1727 881 877 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00864 876 874 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00863 877 875 876 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00862 849 856 852 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00861 1727 848 849 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00860 852 855 851 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00859 1727 851 853 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00858 853 855 850 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00857 850 856 857 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00856 855 856 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00855 1727 1810 856 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00854 857 854 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00853 1727 889 854 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00852 848 852 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00851 1727 852 848 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00850 851 850 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00849 863 862 875 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00848 875 861 863 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00847 863 860 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00846 859 995 858 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00845 1727 859 860 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00844 858 1086 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00843 1727 847 845 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00842 847 969 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00841 1727 844 846 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00840 844 843 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00839 1727 842 841 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00838 842 864 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00837 1727 840 839 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00836 840 980 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00835 1727 819 915 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00834 828 827 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00833 827 830 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00832 1727 762 827 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00831 765 912 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00830 764 1758 834 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00829 1727 765 764 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00828 1727 830 743 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00827 743 829 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00826 907 833 743 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00825 743 834 907 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00824 1727 1758 726 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00823 726 1239 727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00822 727 761 823 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00821 723 819 820 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00820 820 829 723 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00819 723 818 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00818 1727 908 735 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00817 735 828 734 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00816 734 824 818 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00815 829 815 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00814 815 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00813 1727 761 815 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00812 732 1239 824 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00811 824 829 732 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00810 732 823 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00809 1727 759 710 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00808 710 878 705 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00807 705 833 758 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00806 793 791 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00805 1727 1708 791 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00804 699 915 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00803 791 878 699 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00802 1727 794 702 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00801 702 798 809 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00800 809 793 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00799 797 758 757 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00798 1727 797 798 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00797 757 908 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00796 712 803 806 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00795 1727 801 712 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00794 806 802 807 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00793 1727 807 714 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00792 714 802 804 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00791 804 803 715 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00790 802 803 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00789 1727 1810 803 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00788 715 812 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00787 1727 809 812 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00786 801 806 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00785 1727 806 801 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00784 807 804 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00783 1727 1003 751 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00782 751 750 778 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00781 788 787 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00780 787 881 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00779 1727 915 787 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00778 1727 780 861 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00777 861 778 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00776 861 779 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00775 692 801 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00774 1727 1243 692 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00773 692 1244 784 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00772 784 1786 692 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00771 1727 784 785 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00770 1727 1239 752 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00769 752 1169 780 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00768 663 767 768 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00767 1727 843 663 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00766 768 766 771 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00765 1727 771 669 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00764 669 766 770 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00763 770 767 668 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00762 766 767 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00761 1727 1810 767 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00760 668 774 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00759 1727 785 774 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00758 843 768 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00757 1727 768 843 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00756 771 770 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00755 1727 965 750 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00754 1727 1245 736 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00753 736 1245 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00752 1727 737 762 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00751 737 736 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00750 748 912 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00749 1727 1245 745 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00748 749 745 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00747 746 748 749 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00746 747 1245 746 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00745 1727 912 747 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00744 740 739 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00743 1727 1708 739 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00742 738 915 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00741 739 762 738 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00740 744 833 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00739 742 746 741 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00738 1727 744 742 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00737 1727 713 890 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00736 713 730 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00735 733 736 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00734 733 730 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00733 1727 1018 733 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00732 1727 733 731 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00731 1727 995 711 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00730 717 725 716 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00729 1727 1018 717 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00728 716 724 718 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00727 1727 718 720 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00726 720 724 722 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00725 722 725 721 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00724 724 725 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00723 1727 1810 725 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00722 721 719 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00721 1727 820 719 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00720 1018 716 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00719 1727 716 1018 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00718 718 722 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00717 1727 893 730 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00716 830 729 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00715 729 1173 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00714 1727 728 729 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00713 689 711 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00712 691 693 690 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00711 1727 689 691 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00710 709 706 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00709 709 707 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00708 1727 1173 709 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00707 1727 709 708 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00706 703 878 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00705 704 708 794 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00704 1727 703 704 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00703 1727 707 759 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00702 693 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00701 1727 759 693 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00700 1727 698 874 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00699 696 694 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00698 697 695 696 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00697 698 701 697 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00696 679 680 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00695 1727 788 680 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00694 677 683 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00693 680 690 677 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00692 701 700 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00691 700 759 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00690 1727 890 700 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00689 1727 1245 688 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00688 688 761 686 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00687 686 890 687 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00686 687 685 779 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00685 862 1003 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00684 1727 890 862 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00683 684 862 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00682 684 681 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00681 1727 682 684 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00680 1727 684 683 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00679 661 672 660 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00678 1727 995 661 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00677 660 671 662 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00676 1727 662 665 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00675 665 671 666 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00674 666 672 667 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00673 671 672 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00672 1727 1810 672 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00671 667 664 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00670 1727 673 664 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00669 995 660 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00668 1727 660 995 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00667 662 666 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00666 1727 679 676 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00665 676 675 673 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00664 673 670 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00663 1727 1758 678 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00662 678 788 674 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00661 674 995 675 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00660 1727 624 626 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00659 547 623 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00658 548 833 547 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00657 624 1245 548 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00656 1727 741 552 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00655 552 628 635 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00654 635 740 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00653 556 639 631 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00652 1727 1245 556 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00651 631 638 632 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00650 1727 632 558 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00649 558 638 634 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00648 634 639 563 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00647 638 639 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00646 1727 1810 639 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00645 563 637 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00644 1727 635 637 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00643 1245 631 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00642 1727 631 1245 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00641 632 634 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00640 628 626 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00639 1727 625 628 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00638 1727 908 543 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00637 543 622 625 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00636 540 1325 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00635 1727 1244 540 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00634 540 1243 621 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00633 621 618 540 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00632 1727 621 617 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00631 1727 1018 761 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00630 1727 1239 544 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00629 544 761 623 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00628 614 618 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00627 1727 611 614 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00626 1727 890 614 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00625 614 612 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00624 610 614 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00623 530 1201 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00622 1727 1244 530 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00621 530 1243 609 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00620 609 612 530 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00619 1727 609 606 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00618 1727 601 520 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00617 520 1086 707 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00616 706 995 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00615 1727 602 706 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00614 1727 1003 706 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00613 706 610 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00612 598 1003 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00611 1727 602 598 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00610 1727 596 598 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00609 598 610 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00608 1727 1169 515 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00607 515 598 694 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00606 513 1115 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00605 1727 1244 513 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00604 513 1243 590 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00603 590 588 513 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00602 1727 590 587 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00601 592 595 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00600 592 681 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00599 1727 890 592 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00598 1727 592 695 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00597 681 585 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00596 585 995 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00595 1727 596 585 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00594 586 595 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00593 586 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00592 1727 601 586 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00591 1727 586 582 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00590 1727 1169 577 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00589 601 577 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00588 1727 578 601 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00587 1727 1245 497 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00586 497 761 580 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00585 1727 685 493 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00584 493 576 494 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00583 494 1239 492 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00582 492 750 578 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00581 1727 580 576 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00580 574 1007 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00579 1727 750 574 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00578 480 572 566 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00577 1727 564 480 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00576 566 573 567 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00575 1727 567 486 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00574 486 573 571 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00573 571 572 485 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00572 573 572 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00571 1727 1810 572 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00570 485 569 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00569 1727 606 569 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00568 564 566 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00567 1727 566 564 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00566 567 571 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00565 1727 1007 685 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00564 555 557 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00563 555 553 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00562 1727 560 555 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00561 1727 555 554 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00560 562 559 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00559 562 618 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00558 1727 560 562 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00557 1727 562 561 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00556 559 612 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00555 1727 611 559 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00554 551 550 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00553 550 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00552 1727 549 550 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00551 1727 546 549 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00550 546 731 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00549 1727 559 557 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00548 523 612 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00547 1727 521 523 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00546 1727 878 523 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00545 523 602 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00544 1727 522 525 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00543 525 526 524 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00542 524 523 622 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00541 545 965 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00540 1727 728 545 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00539 1727 1007 545 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00538 545 551 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00537 560 545 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00536 1727 1173 833 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00535 529 711 528 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00534 1727 595 531 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00533 528 553 527 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00532 531 588 529 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00531 1727 527 526 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00530 535 542 534 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00529 1727 532 535 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00528 534 541 533 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00527 1727 533 537 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00526 537 541 538 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00525 538 542 539 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00524 541 542 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00523 1727 1810 542 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00522 539 536 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00521 1727 617 536 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00520 532 534 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00519 1727 534 532 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00518 533 538 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00517 516 878 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00516 516 995 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00515 1727 1173 516 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00514 1727 516 514 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00513 510 995 509 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00512 1727 819 511 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00511 509 1086 512 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00510 511 801 510 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00509 1727 512 508 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00508 1727 1086 517 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00507 517 1169 519 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00506 1727 833 518 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00505 522 518 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00504 1727 519 522 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00503 1727 1758 496 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00502 496 506 495 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00501 495 1003 502 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00500 501 500 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00499 1727 506 500 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00498 499 582 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00497 500 498 499 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00496 498 491 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00495 491 682 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00494 1727 1003 491 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00493 505 1173 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00492 507 508 506 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00491 1727 505 507 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00490 1727 501 504 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00489 504 502 503 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00488 503 670 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00487 487 574 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00486 1727 580 487 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00485 1727 488 487 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00484 487 728 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00483 484 487 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00482 1727 478 476 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00481 478 532 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00480 490 488 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00479 1727 728 490 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00478 1727 965 490 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00477 490 489 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00476 682 490 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00475 1727 477 479 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00474 477 848 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00473 481 596 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00472 483 484 482 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00471 1727 481 483 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00470 1727 440 359 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00469 359 439 438 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00468 438 670 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00467 446 448 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00466 1727 445 448 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00465 372 561 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00464 448 444 372 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00463 1727 1758 364 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00462 364 445 360 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00461 360 612 439 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00460 353 434 430 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00459 1727 612 353 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00458 430 436 431 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00457 1727 431 354 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00456 354 436 433 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00455 433 434 355 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00454 436 434 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00453 1727 1810 434 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00452 355 435 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00451 1727 438 435 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00450 612 430 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00449 1727 430 612 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00448 431 433 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00447 440 443 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00446 1727 445 443 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00445 366 554 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00444 443 441 366 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00443 1727 1758 370 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00442 370 521 371 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00441 371 618 444 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00440 1727 618 553 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00439 427 731 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00438 427 965 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00437 1727 1007 427 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00436 1727 427 424 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00435 421 422 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00434 422 622 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00433 1727 915 422 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00432 1727 1086 342 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00431 342 595 420 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00430 1727 1015 335 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00429 335 801 334 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00428 334 711 414 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00427 1727 801 878 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00426 419 417 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00425 419 1173 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00424 1727 420 419 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00423 1727 419 415 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00422 1727 1015 336 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00421 336 801 332 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00420 332 711 417 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00419 1727 1086 596 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00418 402 403 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00417 403 400 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00416 1727 415 403 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00415 327 413 406 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00414 1727 1003 327 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00413 406 412 407 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00412 1727 407 329 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00411 329 412 409 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00410 409 413 330 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00409 412 413 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00408 1727 1810 413 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00407 330 411 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00406 1727 503 411 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00405 1003 406 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00404 1727 406 1003 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00403 407 409 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00402 1727 1086 321 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00401 321 1173 398 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00400 304 381 374 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00399 1727 1086 304 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00398 374 382 373 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00397 1727 373 306 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00396 306 382 377 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00395 377 381 307 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00394 382 381 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00393 1727 1810 381 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00392 307 376 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00391 1727 396 376 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00390 1086 374 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00389 1727 374 1086 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00388 373 377 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00387 1727 395 320 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00386 320 399 396 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00385 396 391 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 1727 401 399 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00383 324 398 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 323 908 324 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 401 402 323 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 1727 965 310 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00379 310 384 380 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00378 1727 576 316 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00377 316 1007 386 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00376 1727 386 385 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00375 384 385 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00374 1727 1708 384 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00373 395 393 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00372 1727 1173 393 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00371 318 482 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00370 393 392 318 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00369 390 488 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00368 1727 386 390 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00367 1727 1086 390 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00366 390 728 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00365 392 390 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00364 1727 446 362 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00363 362 361 363 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00362 363 670 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00361 293 298 365 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00360 1727 618 293 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00359 365 297 368 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00358 1727 368 369 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00357 369 297 367 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00356 367 298 299 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00355 297 298 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00354 1727 1810 298 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00353 299 296 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00352 1727 363 296 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00351 618 365 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00350 1727 365 618 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00349 368 367 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00348 445 356 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00347 356 333 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00346 1727 915 356 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00345 1727 1758 358 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00344 358 445 357 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00343 357 618 361 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00342 1727 612 350 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00341 1727 345 346 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00340 345 424 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00339 1727 595 338 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00338 338 351 340 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00337 340 1086 339 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00336 339 337 341 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00335 349 611 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00334 349 612 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00333 1727 618 349 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00332 1727 349 351 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00331 1727 350 352 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00330 352 893 348 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00329 348 553 347 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00328 343 415 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00327 1727 488 343 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00326 1727 351 343 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00325 343 346 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00324 344 343 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00323 328 347 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00322 328 965 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00321 1727 279 328 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00320 1727 328 400 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00319 1727 1086 281 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00318 281 595 282 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00317 1727 1003 595 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00316 1727 588 277 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00315 277 685 279 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00314 331 282 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00313 1727 414 331 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00312 1727 1173 331 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00311 331 488 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00310 333 331 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00309 391 322 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00308 1727 1708 322 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00307 273 915 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00306 322 596 273 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00305 267 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00304 1727 685 267 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00303 325 488 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00302 325 400 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00301 1727 415 325 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00300 1727 325 326 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00299 253 259 301 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00298 1727 300 253 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00297 301 258 303 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00296 1727 303 305 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00295 305 258 302 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00294 302 259 257 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00293 258 259 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00292 1727 1810 259 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00291 257 256 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00290 1727 587 256 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00289 300 301 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00288 1727 301 300 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00287 303 302 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00286 317 1173 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00285 1727 915 317 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00284 1727 596 317 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00283 317 272 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00282 319 317 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 1727 268 272 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 1727 1758 314 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00279 314 319 311 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 311 965 312 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 309 308 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 1727 319 308 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00275 261 380 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00274 308 315 261 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00273 1727 576 264 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00272 264 1758 265 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00271 313 685 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00270 313 265 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00269 1727 965 313 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00268 1727 313 315 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 233 234 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00266 1727 1708 234 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00265 180 915 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00264 234 611 180 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00263 1727 588 611 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 240 238 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00261 240 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00260 1727 350 240 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00259 1727 240 441 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00258 237 236 181 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00257 1727 237 238 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00256 181 588 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00255 182 250 247 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00254 1727 819 182 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00253 247 252 244 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00252 1727 244 183 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00251 183 252 246 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00250 246 250 185 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00249 252 250 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00248 1727 1810 250 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00247 185 251 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00246 1727 248 251 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00245 819 247 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 1727 247 819 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 244 246 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00242 1727 231 521 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00241 231 230 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00240 236 553 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00239 1727 230 236 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00238 1727 229 230 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 229 728 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00236 1727 424 229 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00235 1727 227 337 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 227 229 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00233 179 488 226 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 226 341 179 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 179 1015 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 1727 224 670 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 223 1003 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00228 1727 521 223 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00227 1727 596 223 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00226 223 1015 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00225 216 217 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00224 1727 514 217 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00223 177 226 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00222 217 219 177 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00221 1727 1169 178 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 178 223 219 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 214 215 176 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 1727 214 213 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 176 1007 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 215 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00215 1727 576 215 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00214 1727 204 202 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 1727 213 173 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00212 173 203 1727 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00211 204 272 174 1727 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00210 174 267 1727 1727 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00209 173 268 204 1727 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00208 206 1239 175 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 1727 206 268 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 175 1169 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00205 212 965 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00204 1727 215 212 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00203 1727 596 212 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00202 212 728 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00201 1727 489 203 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 489 201 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 201 265 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00198 1727 1007 201 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00197 1727 187 186 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 187 300 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00195 1727 309 172 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00194 172 312 198 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00193 198 670 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 169 197 193 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00191 1727 965 169 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00190 193 196 190 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00189 1727 190 170 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00188 170 196 192 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00187 192 197 171 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00186 196 197 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00185 1727 1810 197 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00184 171 194 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00183 1727 198 194 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00182 965 193 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00181 1727 193 965 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 190 192 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00179 162 588 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00178 1727 155 160 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00177 157 160 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 158 162 157 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 159 155 158 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 1727 588 159 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 248 1708 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00172 1727 166 248 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00171 1727 154 155 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 154 236 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00169 137 908 136 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 1727 137 138 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 136 1239 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 1727 819 168 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00165 168 163 166 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00164 166 165 167 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00163 167 184 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 1727 184 163 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00161 165 819 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00160 141 143 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 1727 1708 143 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00158 142 915 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00157 143 728 142 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00156 1727 1015 602 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00155 1727 344 139 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 139 138 146 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00153 146 141 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 1727 421 135 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 135 132 134 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 134 1708 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 144 152 145 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00148 1727 1239 144 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00147 145 153 147 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00146 1727 147 151 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00145 151 153 150 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00144 150 152 148 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00143 153 152 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00142 1727 1810 152 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00141 148 149 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00140 1727 146 149 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00139 1239 145 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 1727 145 1239 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 147 150 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00136 113 121 114 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00135 1727 1015 113 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00134 114 120 115 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00133 1727 115 116 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00132 116 120 118 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00131 118 121 117 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00130 120 121 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00129 1727 1810 121 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00128 117 119 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00127 1727 127 119 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00126 1015 114 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 1727 114 1015 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 115 118 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00123 1727 216 129 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00122 129 125 127 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00121 127 128 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 105 1173 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00119 1727 915 105 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00118 1727 1015 124 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 124 514 125 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 125 122 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 128 131 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 1727 1708 131 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00113 130 915 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00112 131 602 130 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00111 1727 1169 111 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 111 212 112 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 1727 267 99 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00108 102 99 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 1727 105 102 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00106 98 101 97 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00105 97 102 98 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00104 1727 224 97 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00103 96 98 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 1727 104 101 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 106 202 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 107 112 106 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 104 105 107 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00098 108 109 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 1727 1708 109 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00096 110 915 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00095 109 488 110 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00094 1727 1239 728 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 84 92 86 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00092 1727 1007 84 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00091 86 91 85 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00090 1727 85 89 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00089 89 91 88 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00088 88 92 90 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00087 91 92 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00086 1727 1810 92 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00085 90 87 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00084 1727 96 87 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00083 1007 86 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 1727 86 1007 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 85 88 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00080 94 576 93 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 1727 94 95 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 93 1239 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 1727 588 15 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 15 333 70 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00075 70 65 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 18 81 78 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00073 1727 588 18 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00072 78 83 75 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00071 1727 75 19 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00070 19 83 77 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 77 81 20 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00068 83 81 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00067 1727 1810 81 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00066 20 82 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00065 1727 79 82 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00064 588 78 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 1727 78 588 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 75 77 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00061 1727 73 16 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 16 70 79 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 79 233 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 1727 908 65 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 72 333 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 17 158 73 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 1727 72 17 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 1727 54 132 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 12 63 56 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00052 1727 54 12 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00051 56 62 57 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00050 1727 57 13 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00049 13 62 59 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00048 59 63 14 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 62 63 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 1727 1810 63 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 14 61 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00044 1727 134 61 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00043 54 56 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 1727 56 54 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 57 59 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00040 1727 819 52 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00039 908 52 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 1727 54 908 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00037 1727 54 11 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 11 819 224 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 1727 1169 488 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 1727 908 122 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 1727 46 45 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 8 326 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 9 48 8 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 46 908 9 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 1727 45 7 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 7 41 42 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 42 108 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 1 33 24 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00025 1727 1169 1 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00024 24 34 28 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 1727 28 3 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 3 34 30 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00021 30 33 2 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 34 33 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00019 1727 1810 33 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 2 32 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 1727 42 32 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 1169 24 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 1727 24 1169 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 28 30 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 1727 1169 10 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 10 1173 48 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 37 95 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 1727 1169 35 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 4 35 1727 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 39 37 4 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 5 1169 39 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 1727 95 5 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 40 1173 1727 1727 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 6 39 41 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 1727 40 6 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 1727 21 22 1727 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 21 564 1727 1727 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
C1812 21 1727 1.568e-14
C1811 22 1727 2.659e-14
C1809 24 1727 2.871e-14
C1805 28 1727 2.005e-14
C1803 30 1727 2.632e-14
C1801 32 1727 2.321e-14
C1800 33 1727 5.165e-14
C1799 34 1727 4.869e-14
C1798 35 1727 2.596e-14
C1796 37 1727 2.16e-14
C1795 38 1727 9.7e-15
C1794 39 1727 5.34e-14
C1793 40 1727 1.662e-14
C1792 41 1727 5.211e-14
C1791 42 1727 7.508e-14
C1790 43 1727 6.05e-15
C1789 44 1727 6.05e-15
C1788 45 1727 4.875e-14
C1787 46 1727 2.605e-14
C1785 48 1727 4.791e-14
C1781 52 1727 1.677e-14
C1780 53 1727 6.05e-15
C1779 54 1727 1.423e-13
C1777 56 1727 2.871e-14
C1776 57 1727 2.005e-14
C1774 59 1727 2.632e-14
C1772 61 1727 2.321e-14
C1771 62 1727 4.869e-14
C1770 63 1727 5.165e-14
C1769 64 1727 6.05e-15
C1768 65 1727 5.559e-14
C1766 67 1727 6.05e-15
C1763 70 1727 5.227e-14
C1762 71 1727 6.05e-15
C1761 72 1727 1.662e-14
C1760 73 1727 4.821e-14
C1758 75 1727 2.005e-14
C1756 77 1727 2.632e-14
C1755 78 1727 2.871e-14
C1754 79 1727 7.628e-14
C1752 81 1727 5.165e-14
C1751 82 1727 2.321e-14
C1750 83 1727 4.869e-14
C1748 85 1727 2.005e-14
C1747 86 1727 2.871e-14
C1746 87 1727 2.321e-14
C1745 88 1727 2.632e-14
C1742 91 1727 4.869e-14
C1741 92 1727 5.165e-14
C1739 94 1727 1.8635e-14
C1738 95 1727 7.089e-14
C1737 96 1727 6.318e-14
C1736 97 1727 4.11e-15
C1735 98 1727 1.853e-14
C1734 99 1727 1.677e-14
C1732 101 1727 5.265e-14
C1731 102 1727 5.219e-14
C1729 104 1727 2.605e-14
C1728 105 1727 8.819e-14
C1725 108 1727 5.579e-14
C1724 109 1727 1.767e-14
C1721 112 1727 5.751e-14
C1719 114 1727 2.871e-14
C1718 115 1727 2.005e-14
C1715 118 1727 2.632e-14
C1714 119 1727 2.321e-14
C1713 120 1727 4.869e-14
C1712 121 1727 5.165e-14
C1711 122 1727 5.271e-14
C1710 123 1727 6.05e-15
C1708 125 1727 4.747e-14
C1707 126 1727 6.05e-15
C1706 127 1727 5.828e-14
C1705 128 1727 5.507e-14
C1702 131 1727 1.767e-14
C1701 132 1727 5.409e-14
C1700 133 1727 6.05e-15
C1699 134 1727 6.956e-14
C1696 137 1727 1.8635e-14
C1695 138 1727 5.233e-14
C1693 140 1727 6.05e-15
C1692 141 1727 5.747e-14
C1690 143 1727 1.767e-14
C1688 145 1727 2.871e-14
C1687 146 1727 7.268e-14
C1686 147 1727 2.005e-14
C1684 149 1727 2.321e-14
C1683 150 1727 2.632e-14
C1681 152 1727 5.165e-14
C1680 153 1727 4.869e-14
C1679 154 1727 1.568e-14
C1678 155 1727 6.133e-14
C1677 156 1727 9.7e-15
C1675 158 1727 6.06e-14
C1673 160 1727 2.596e-14
C1671 162 1727 2.16e-14
C1670 163 1727 2.596e-14
C1668 164 1727 7.76e-15
C1667 165 1727 2.16e-14
C1666 166 1727 5.454e-14
C1659 173 1727 4.11e-15
C1653 179 1727 4.11e-15
C1648 184 1727 5.024e-14
C1645 186 1727 2.899e-14
C1644 187 1727 1.568e-14
C1641 190 1727 2.005e-14
C1639 192 1727 2.632e-14
C1638 193 1727 2.871e-14
C1637 194 1727 2.321e-14
C1635 196 1727 4.869e-14
C1634 197 1727 5.165e-14
C1633 198 1727 5.108e-14
C1632 199 1727 6.05e-15
C1630 201 1727 1.8635e-14
C1629 202 1727 5.079e-14
C1628 203 1727 4.494e-14
C1627 204 1727 2.299e-14
C1625 206 1727 1.8635e-14
C1624 207 1727 8.58e-15
C1619 212 1727 7.266e-14
C1618 213 1727 6.658e-14
C1617 214 1727 1.8635e-14
C1616 215 1727 8.253e-14
C1615 216 1727 6.527e-14
C1614 217 1727 1.767e-14
C1613 218 1727 6.05e-15
C1612 219 1727 4.817e-14
C1608 223 1727 6.306e-14
C1607 224 1727 1.8722e-13
C1605 226 1727 6.977e-14
C1604 227 1727 1.568e-14
C1602 229 1727 8.616e-14
C1601 230 1727 8.939e-14
C1600 231 1727 1.568e-14
C1598 233 1727 7.427e-14
C1597 234 1727 1.767e-14
C1596 235 1727 6.05e-15
C1595 236 1727 9.192e-14
C1594 237 1727 1.8635e-14
C1593 238 1727 5.203e-14
C1591 240 1727 2.455e-14
C1587 244 1727 2.005e-14
C1585 246 1727 2.632e-14
C1584 247 1727 2.871e-14
C1583 248 1727 5.882e-14
C1581 250 1727 5.165e-14
C1580 251 1727 2.321e-14
C1579 252 1727 4.869e-14
C1575 256 1727 2.321e-14
C1573 258 1727 4.869e-14
C1572 259 1727 5.165e-14
C1571 260 1727 6.05e-15
C1566 265 1727 8.776e-14
C1564 267 1727 1.1581e-13
C1563 268 1727 7.867e-14
C1559 272 1727 7.27e-14
C1555 276 1727 6.05e-15
C1552 279 1727 5.031e-14
C1549 282 1727 5.061e-14
C1539 292 1727 6.05e-15
C1534 296 1727 2.321e-14
C1533 297 1727 4.869e-14
C1532 298 1727 5.165e-14
C1530 300 1727 6.919e-14
C1529 301 1727 2.871e-14
C1528 302 1727 2.632e-14
C1527 303 1727 2.005e-14
C1522 308 1727 1.767e-14
C1521 309 1727 6.407e-14
C1518 312 1727 5.505e-14
C1517 313 1727 2.455e-14
C1515 315 1727 5.323e-14
C1513 317 1727 2.72e-14
C1511 319 1727 1.0481e-13
C1508 322 1727 1.767e-14
C1505 325 1727 2.455e-14
C1504 326 1727 8.027e-14
C1502 328 1727 2.455e-14
C1499 331 1727 2.72e-14
C1497 333 1727 2.2511e-13
C1493 337 1727 7.216e-14
C1489 341 1727 5.561e-14
C1487 343 1727 2.72e-14
C1486 344 1727 7.579e-14
C1485 345 1727 1.568e-14
C1484 346 1727 4.573e-14
C1483 347 1727 9.915e-14
C1481 349 1727 2.455e-14
C1480 350 1727 1.17e-13
C1479 351 1727 1.0673e-13
C1474 356 1727 1.8635e-14
C1469 361 1727 5.625e-14
C1467 363 1727 6.308e-14
C1465 365 1727 2.871e-14
C1463 367 1727 2.632e-14
C1462 368 1727 2.005e-14
C1456 373 1727 2.005e-14
C1455 374 1727 2.871e-14
C1453 376 1727 2.321e-14
C1452 377 1727 2.632e-14
C1449 380 1727 5.331e-14
C1448 381 1727 5.165e-14
C1447 382 1727 4.869e-14
C1445 384 1727 5.568e-14
C1444 385 1727 1.677e-14
C1443 386 1727 8.286e-14
C1439 390 1727 2.72e-14
C1438 391 1727 6.707e-14
C1437 392 1727 5.535e-14
C1436 393 1727 1.767e-14
C1435 394 1727 6.05e-15
C1434 395 1727 5.447e-14
C1433 396 1727 8.228e-14
C1432 397 1727 6.05e-15
C1431 398 1727 4.761e-14
C1430 399 1727 5.265e-14
C1429 400 1727 1.0082e-13
C1428 401 1727 2.605e-14
C1427 402 1727 4.151e-14
C1426 403 1727 1.8635e-14
C1423 406 1727 2.871e-14
C1422 407 1727 2.005e-14
C1420 409 1727 2.632e-14
C1418 411 1727 2.321e-14
C1417 412 1727 4.869e-14
C1416 413 1727 5.165e-14
C1415 414 1727 6.243e-14
C1414 415 1727 1.6737e-13
C1412 417 1727 5.355e-14
C1410 419 1727 2.455e-14
C1409 420 1727 4.551e-14
C1408 421 1727 7.391e-14
C1407 422 1727 1.8635e-14
C1405 424 1727 9.671e-14
C1402 427 1727 2.455e-14
C1399 430 1727 2.871e-14
C1398 431 1727 2.005e-14
C1396 433 1727 2.632e-14
C1395 434 1727 5.165e-14
C1394 435 1727 2.321e-14
C1393 436 1727 4.869e-14
C1392 437 1727 6.05e-15
C1391 438 1727 5.348e-14
C1390 439 1727 5.025e-14
C1389 440 1727 5.567e-14
C1388 441 1727 7.243e-14
C1387 442 1727 6.05e-15
C1386 443 1727 1.767e-14
C1385 444 1727 5.591e-14
C1384 445 1727 1.8134e-13
C1383 446 1727 6.887e-14
C1382 447 1727 6.05e-15
C1381 448 1727 1.767e-14
C1373 456 1727 6.05e-15
C1372 457 1727 6.05e-15
C1352 476 1727 5.803e-14
C1351 477 1727 1.568e-14
C1350 478 1727 1.568e-14
C1349 479 1727 2.899e-14
C1347 481 1727 1.662e-14
C1346 482 1727 9.051e-14
C1344 484 1727 5.454e-14
C1341 487 1727 2.72e-14
C1340 488 1727 3.9774e-13
C1339 489 1727 1.094e-13
C1338 490 1727 2.72e-14
C1337 491 1727 1.8635e-14
C1330 498 1727 5.947e-14
C1328 500 1727 1.767e-14
C1327 501 1727 5.447e-14
C1326 502 1727 6.225e-14
C1325 503 1727 8.348e-14
C1323 505 1727 1.662e-14
C1322 506 1727 9.403e-14
C1320 508 1727 5.75e-14
C1316 512 1727 2.306e-14
C1315 513 1727 7.43e-15
C1314 514 1727 1.2938e-13
C1312 516 1727 2.455e-14
C1310 518 1727 1.677e-14
C1309 519 1727 5.346e-14
C1307 521 1727 2.4568e-13
C1306 522 1727 6.753e-14
C1305 523 1727 5.596e-14
C1302 526 1727 5.62e-14
C1301 527 1727 2.306e-14
C1298 530 1727 7.43e-15
C1296 532 1727 2.0599e-13
C1295 533 1727 2.005e-14
C1294 534 1727 2.871e-14
C1292 536 1727 2.321e-14
C1290 538 1727 2.632e-14
C1288 540 1727 7.43e-15
C1287 541 1727 4.869e-14
C1286 542 1727 5.165e-14
C1283 545 1727 2.72e-14
C1282 546 1727 1.568e-14
C1279 549 1727 5.053e-14
C1278 550 1727 1.8635e-14
C1277 551 1727 5.321e-14
C1275 553 1727 2.5674e-13
C1274 554 1727 5.597e-14
C1273 555 1727 2.455e-14
C1271 557 1727 4.419e-14
C1269 559 1727 9.582e-14
C1268 560 1727 1.1978e-13
C1267 561 1727 5.837e-14
C1266 562 1727 2.455e-14
C1263 564 1727 1.3207e-13
C1261 566 1727 2.871e-14
C1260 567 1727 2.005e-14
C1258 569 1727 2.321e-14
C1256 571 1727 2.632e-14
C1255 572 1727 5.165e-14
C1254 573 1727 4.869e-14
C1253 574 1727 6.091e-14
C1251 576 1727 2.6485e-13
C1250 577 1727 1.677e-14
C1249 578 1727 5.816e-14
C1247 580 1727 1.04e-13
C1245 582 1727 5.717e-14
C1242 585 1727 1.8635e-14
C1241 586 1727 2.455e-14
C1240 587 1727 1.289e-13
C1239 588 1727 4.967e-13
C1237 590 1727 2.639e-14
C1235 592 1727 2.455e-14
C1232 595 1727 2.8916e-13
C1231 596 1727 3.9774e-13
C1229 598 1727 6.306e-14
C1226 601 1727 1.2784e-13
C1225 602 1727 1.9067e-13
C1221 606 1727 1.5626e-13
C1218 609 1727 2.639e-14
C1217 610 1727 1.052e-13
C1216 611 1727 2.5235e-13
C1215 612 1727 3.5332e-13
C1213 614 1727 2.72e-14
C1210 617 1727 5.834e-14
C1209 618 1727 3.4465e-13
C1206 621 1727 2.639e-14
C1205 622 1727 1.4535e-13
C1204 623 1727 5.001e-14
C1203 624 1727 2.605e-14
C1202 625 1727 6.696e-14
C1201 626 1727 5.85e-14
C1199 628 1727 5.041e-14
C1198 629 1727 6.05e-15
C1196 631 1727 2.871e-14
C1195 632 1727 2.005e-14
C1193 634 1727 2.632e-14
C1192 635 1727 6.308e-14
C1190 637 1727 2.321e-14
C1189 638 1727 4.869e-14
C1188 639 1727 5.165e-14
C1184 643 1727 6.05e-15
C1183 644 1727 6.05e-15
C1169 658 1727 6.05e-15
C1167 659 1727 9.7e-15
C1166 660 1727 2.871e-14
C1164 662 1727 2.005e-14
C1162 664 1727 2.321e-14
C1160 666 1727 2.632e-14
C1156 670 1727 4.4587e-13
C1155 671 1727 4.869e-14
C1154 672 1727 5.165e-14
C1153 673 1727 5.108e-14
C1151 675 1727 4.785e-14
C1147 679 1727 5.087e-14
C1146 680 1727 1.767e-14
C1145 681 1727 1.1238e-13
C1144 682 1727 1.1174e-13
C1143 683 1727 4.637e-14
C1142 684 1727 2.455e-14
C1141 685 1727 2.4807e-13
C1137 689 1727 1.662e-14
C1136 690 1727 6.737e-14
C1134 692 1727 7.43e-15
C1133 693 1727 5.766e-14
C1132 694 1727 5.481e-14
C1131 695 1727 5.897e-14
C1128 698 1727 2.605e-14
C1126 700 1727 1.8635e-14
C1125 701 1727 4.151e-14
C1123 703 1727 1.662e-14
C1120 706 1727 5.431e-14
C1119 707 1727 8.61e-14
C1118 708 1727 6.322e-14
C1117 709 1727 2.455e-14
C1115 711 1727 2.3819e-13
C1113 713 1727 1.568e-14
C1110 716 1727 2.871e-14
C1108 718 1727 2.005e-14
C1107 719 1727 2.321e-14
C1104 722 1727 2.632e-14
C1103 723 1727 4.11e-15
C1102 724 1727 4.869e-14
C1101 725 1727 5.165e-14
C1098 728 1727 4.8822e-13
C1097 729 1727 1.8635e-14
C1096 730 1727 1.1954e-13
C1095 731 1727 1.3988e-13
C1094 732 1727 4.11e-15
C1093 733 1727 2.455e-14
C1090 736 1727 8.448e-14
C1089 737 1727 1.568e-14
C1087 739 1727 1.767e-14
C1086 740 1727 5.747e-14
C1085 741 1727 5.781e-14
C1083 743 1727 7.43e-15
C1082 744 1727 1.662e-14
C1081 745 1727 2.596e-14
C1080 746 1727 6.06e-14
C1078 748 1727 2.16e-14
C1076 750 1727 1.2364e-13
C1070 756 1727 6.05e-15
C1068 758 1727 4.571e-14
C1067 759 1727 1.387e-13
C1065 761 1727 3.1771e-13
C1064 762 1727 8.068e-14
C1061 765 1727 1.662e-14
C1059 766 1727 4.869e-14
C1058 767 1727 5.165e-14
C1057 768 1727 2.871e-14
C1055 770 1727 2.632e-14
C1054 771 1727 2.005e-14
C1051 774 1727 2.321e-14
C1047 778 1727 5.991e-14
C1046 779 1727 6.026e-14
C1045 780 1727 5.106e-14
C1041 784 1727 2.639e-14
C1040 785 1727 8.114e-14
C1038 787 1727 1.8635e-14
C1037 788 1727 1.1781e-13
C1034 791 1727 1.767e-14
C1033 792 1727 6.05e-15
C1032 793 1727 5.987e-14
C1031 794 1727 5.061e-14
C1030 795 1727 6.05e-15
C1028 797 1727 1.8635e-14
C1027 798 1727 4.633e-14
C1026 799 1727 6.05e-15
C1025 800 1727 6.05e-15
C1024 801 1727 3.0672e-13
C1023 802 1727 4.869e-14
C1022 803 1727 5.165e-14
C1021 804 1727 2.632e-14
C1019 806 1727 2.871e-14
C1018 807 1727 2.005e-14
C1017 808 1727 6.05e-15
C1016 809 1727 7.988e-14
C1013 812 1727 2.321e-14
C1010 815 1727 1.8635e-14
C1007 818 1727 7.575e-14
C1006 819 1727 5.8602e-13
C1005 820 1727 5.298e-14
C1002 823 1727 5.895e-14
C1001 824 1727 5.192e-14
C999 826 1727 6.05e-15
C998 827 1727 1.8635e-14
C997 828 1727 5.496e-14
C996 829 1727 1.4158e-13
C995 830 1727 1.1631e-13
C992 833 1727 3.3716e-13
C991 834 1727 4.821e-14
C985 839 1727 9.235e-14
C984 840 1727 1.568e-14
C983 841 1727 6.643e-14
C982 842 1727 1.568e-14
C981 843 1727 7.687e-14
C980 844 1727 1.568e-14
C979 845 1727 5.875e-14
C978 846 1727 3.907e-14
C977 847 1727 1.568e-14
C976 848 1727 1.2007e-13
C974 850 1727 2.632e-14
C973 851 1727 2.005e-14
C972 852 1727 2.871e-14
C970 854 1727 2.321e-14
C969 855 1727 4.869e-14
C968 856 1727 5.165e-14
C965 859 1727 1.8635e-14
C964 860 1727 5.263e-14
C963 861 1727 5.209e-14
C962 862 1727 8.71e-14
C961 863 1727 4.11e-15
C960 864 1727 1.1167e-13
C958 866 1727 2.871e-14
C957 867 1727 2.005e-14
C956 868 1727 2.321e-14
C954 870 1727 2.632e-14
C952 872 1727 4.869e-14
C951 873 1727 5.165e-14
C950 874 1727 6.825e-14
C949 875 1727 6.943e-14
C947 877 1727 1.767e-14
C946 878 1727 2.7006e-13
C945 879 1727 1.8635e-14
C944 880 1727 5.319e-14
C943 881 1727 1.3443e-13
C941 883 1727 7.607e-14
C940 884 1727 4.747e-14
C939 885 1727 1.767e-14
C937 887 1727 5.507e-14
C935 889 1727 1.361e-13
C934 890 1727 3.0438e-13
C933 891 1727 2.639e-14
C932 892 1727 7.43e-15
C931 893 1727 2.6587e-13
C929 895 1727 2.871e-14
C927 897 1727 2.005e-14
C926 898 1727 8.348e-14
C925 899 1727 2.321e-14
C924 900 1727 2.632e-14
C922 902 1727 4.869e-14
C921 903 1727 5.165e-14
C919 905 1727 2.605e-14
C917 907 1727 7.457e-14
C916 908 1727 6.2046e-13
C915 909 1727 6.221e-14
C913 911 1727 1.767e-14
C912 912 1727 1.3662e-13
C910 914 1727 1.8635e-14
C909 915 1727 7.95029e-13
C908 916 1727 1.677e-14
C905 919 1727 2.632e-14
C904 920 1727 2.871e-14
C903 921 1727 2.005e-14
C901 923 1727 2.321e-14
C900 924 1727 4.869e-14
C899 925 1727 5.165e-14
C895 929 1727 7.43e-15
C888 936 1727 7.43e-15
C887 937 1727 7.43e-15
C886 938 1727 7.43e-15
C885 939 1727 7.43e-15
C884 940 1727 7.43e-15
C877 947 1727 7.43e-15
C875 948 1727 1.568e-14
C874 949 1727 2.539e-14
C873 950 1727 6.727e-14
C871 952 1727 2.005e-14
C869 954 1727 2.632e-14
C868 955 1727 2.871e-14
C866 957 1727 2.321e-14
C864 959 1727 4.869e-14
C861 962 1727 4.994e-14
C860 963 1727 5.165e-14
C858 965 1727 5.9558e-13
C857 966 1727 2.639e-14
C854 969 1727 9.247e-14
C852 971 1727 2.005e-14
C851 972 1727 2.871e-14
C848 975 1727 2.321e-14
C846 977 1727 2.632e-14
C845 978 1727 4.869e-14
C843 980 1727 1.3303e-13
C842 981 1727 5.165e-14
C838 985 1727 2.871e-14
C837 986 1727 2.005e-14
C835 988 1727 4.869e-14
C834 989 1727 2.321e-14
C832 991 1727 2.632e-14
C831 992 1727 5.165e-14
C830 993 1727 7.514e-14
C828 995 1727 4.8135e-13
C826 997 1727 2.639e-14
C822 1001 1727 7.802e-14
C820 1003 1727 5.1506e-13
C819 1004 1727 2.639e-14
C816 1007 1727 6.0754e-13
C813 1010 1727 2.639e-14
C812 1011 1727 8.58e-15
C811 1012 1727 8.594e-14
C808 1015 1727 4.022e-13
C807 1016 1727 2.639e-14
C805 1018 1727 2.4756e-13
C804 1019 1727 2.639e-14
C802 1021 1727 7.43e-15
C799 1024 1727 2.871e-14
C798 1025 1727 9.7e-15
C797 1026 1727 2.005e-14
C796 1027 1727 7.158e-14
C794 1029 1727 2.632e-14
C792 1031 1727 5.165e-14
C791 1032 1727 2.321e-14
C790 1033 1727 4.869e-14
C787 1036 1727 1.8635e-14
C781 1042 1727 7.71e-14
C780 1043 1727 4.696e-14
C779 1044 1727 7.939e-14
C778 1045 1727 7.79e-15
C776 1047 1727 6.256e-14
C775 1048 1727 7.43e-15
C774 1049 1727 2.9265e-14
C773 1050 1727 1.1098e-13
C771 1052 1727 5.087e-14
C766 1057 1727 4.849e-14
C765 1058 1727 2.72e-14
C761 1061 1727 2.371e-14
C760 1062 1727 1.568e-14
C759 1063 1727 1.568e-14
C758 1064 1727 7.207e-14
C756 1066 1727 2.871e-14
C755 1067 1727 2.005e-14
C752 1070 1727 2.632e-14
C751 1071 1727 4.869e-14
C750 1072 1727 5.165e-14
C749 1073 1727 2.321e-14
C747 1075 1727 8.887e-14
C746 1076 1727 2.871e-14
C745 1077 1727 1.3274e-13
C744 1078 1727 2.005e-14
C743 1079 1727 2.321e-14
C742 1080 1727 2.632e-14
C739 1083 1727 4.869e-14
C738 1084 1727 5.165e-14
C737 1085 1727 7.154e-14
C736 1086 1727 6.1761e-13
C735 1087 1727 2.639e-14
C734 1088 1727 7.43e-15
C732 1090 1727 1.662e-14
C730 1092 1727 2.871e-14
C729 1093 1727 2.005e-14
C727 1095 1727 2.632e-14
C725 1097 1727 4.869e-14
C724 1098 1727 5.165e-14
C723 1099 1727 2.321e-14
C722 1100 1727 5.29e-14
C721 1101 1727 4.11e-15
C719 1103 1727 2.299e-14
C718 1104 1727 7.817e-14
C716 1106 1727 2.445e-14
C714 1108 1727 2.596e-14
C712 1110 1727 5.365e-14
C710 1112 1727 2.16e-14
C709 1113 1727 1.568e-14
C708 1114 1727 5.409e-14
C707 1115 1727 2.8864e-13
C705 1117 1727 2.005e-14
C704 1118 1727 2.871e-14
C703 1119 1727 2.632e-14
C700 1122 1727 9.074e-14
C699 1123 1727 2.321e-14
C698 1124 1727 4.869e-14
C697 1125 1727 5.165e-14
C695 1127 1727 6.066e-14
C694 1128 1727 5.386e-14
C693 1129 1727 5.516e-14
C689 1133 1727 6.052e-14
C688 1134 1727 5.826e-14
C683 1139 1727 7.43e-15
C682 1140 1727 7.43e-15
C665 1156 1727 1.568e-14
C664 1157 1727 2.371e-14
C661 1160 1727 2.005e-14
C659 1162 1727 2.871e-14
C658 1163 1727 4.869e-14
C657 1164 1727 2.321e-14
C656 1165 1727 2.632e-14
C654 1167 1727 5.234e-14
C653 1168 1727 5.165e-14
C652 1169 1727 6.7571e-13
C650 1171 1727 2.639e-14
C648 1173 1727 9.16849e-13
C645 1176 1727 2.639e-14
C644 1177 1727 8.31e-14
C643 1178 1727 5.874e-14
C638 1183 1727 9.7e-15
C637 1184 1727 2.596e-14
C636 1185 1727 6.597e-14
C635 1186 1727 2.16e-14
C634 1187 1727 5.986e-14
C633 1188 1727 4.881e-14
C632 1189 1727 1.8635e-14
C631 1190 1727 1.6207e-13
C629 1192 1727 2.871e-14
C628 1193 1727 7.154e-14
C627 1194 1727 2.005e-14
C625 1196 1727 2.632e-14
C623 1198 1727 5.165e-14
C622 1199 1727 4.869e-14
C621 1200 1727 2.321e-14
C620 1201 1727 2.9986e-13
C619 1202 1727 6.286e-14
C618 1203 1727 1.8635e-14
C617 1204 1727 8.611e-14
C615 1206 1727 2.0171e-13
C614 1207 1727 8.736e-14
C613 1208 1727 4.959e-14
C612 1209 1727 2.605e-14
C610 1211 1727 1.8635e-14
C608 1213 1727 2.871e-14
C607 1214 1727 2.005e-14
C605 1216 1727 2.632e-14
C603 1218 1727 2.321e-14
C602 1219 1727 5.165e-14
C601 1220 1727 4.869e-14
C600 1221 1727 5.598e-14
C599 1222 1727 1.767e-14
C598 1223 1727 6.05e-15
C597 1224 1727 5.981e-14
C596 1225 1727 1.3866e-13
C595 1226 1727 4.839e-14
C594 1227 1727 2.605e-14
C593 1228 1727 2.371e-14
C592 1229 1727 7.567e-14
C587 1234 1727 2.321e-14
C586 1235 1727 4.869e-14
C583 1238 1727 5.165e-14
C582 1239 1727 7.9007e-13
C580 1241 1727 6.074e-14
C579 1242 1727 7.43e-15
C578 1243 1727 6.5656e-13
C577 1244 1727 7.7518e-13
C576 1245 1727 4.8735e-13
C575 1246 1727 7.43e-15
C572 1249 1727 7.76e-15
C568 1253 1727 4.11e-15
C564 1257 1727 6.138e-14
C562 1259 1727 4.869e-14
C561 1260 1727 2.321e-14
C557 1264 1727 5.165e-14
C556 1265 1727 1.0802e-13
C554 1267 1727 1.0521e-13
C550 1271 1727 5.291e-14
C545 1276 1727 4.981e-14
C540 1281 1727 5.647e-14
C539 1282 1727 1.0275e-13
C536 1285 1727 4.11e-15
C535 1286 1727 7.577e-14
C533 1288 1727 6.636e-14
C528 1293 1727 8.587e-14
C525 1295 1727 1.568e-14
C524 1296 1727 2.871e-14
C523 1297 1727 2.005e-14
C522 1298 1727 2.632e-14
C520 1300 1727 2.639e-14
C517 1303 1727 2.445e-14
C514 1306 1727 2.596e-14
C513 1307 1727 2.16e-14
C512 1308 1727 1.6881e-13
C510 1310 1727 4.929e-14
C509 1311 1727 2.871e-14
C507 1313 1727 2.005e-14
C506 1314 1727 2.632e-14
C504 1316 1727 4.11e-15
C503 1317 1727 2.455e-14
C501 1319 1727 1.8635e-14
C499 1321 1727 7.43e-15
C498 1322 1727 2.72e-14
C495 1325 1727 3.8066e-13
C494 1326 1727 4.7267e-13
C491 1329 1727 2.605e-14
C487 1333 1727 1.0266e-13
C486 1334 1727 4.103e-14
C483 1337 1727 4.581e-14
C482 1338 1727 8.505e-14
C481 1339 1727 2.72e-14
C479 1341 1727 1.8635e-14
C475 1344 1727 6.919e-14
C474 1345 1727 3.067e-14
C473 1346 1727 1.568e-14
C472 1347 1727 1.568e-14
C471 1348 1727 1.568e-14
C470 1349 1727 6.727e-14
C469 1350 1727 2.005e-14
C468 1351 1727 2.871e-14
C466 1353 1727 5.114e-14
C465 1354 1727 2.321e-14
C463 1356 1727 2.632e-14
C462 1357 1727 4.869e-14
C460 1359 1727 9.847e-14
C459 1360 1727 5.165e-14
C458 1361 1727 2.005e-14
C456 1363 1727 2.871e-14
C454 1365 1727 6.794e-14
C453 1366 1727 2.321e-14
C451 1368 1727 2.632e-14
C450 1369 1727 4.869e-14
C449 1370 1727 5.867e-14
C448 1371 1727 5.165e-14
C445 1374 1727 2.455e-14
C444 1375 1727 5.181e-14
C443 1376 1727 7.95e-14
C442 1377 1727 1.8635e-14
C440 1379 1727 1.662e-14
C439 1380 1727 8.142e-14
C437 1382 1727 5.541e-14
C435 1384 1727 5.293e-14
C434 1385 1727 6.05e-15
C433 1386 1727 1.767e-14
C432 1387 1727 2.005e-14
C431 1388 1727 2.871e-14
C429 1390 1727 6.798e-14
C428 1391 1727 2.321e-14
C425 1394 1727 2.632e-14
C424 1395 1727 4.869e-14
C423 1396 1727 5.165e-14
C419 1400 1727 5.221e-14
C418 1401 1727 7.43e-15
C417 1402 1727 2.445e-14
C416 1403 1727 4.951e-14
C414 1405 1727 7.631e-14
C413 1406 1727 7.994e-14
C411 1408 1727 1.8635e-14
C410 1409 1727 1.0535e-13
C409 1410 1727 2.0045e-13
C407 1412 1727 2.455e-14
C405 1414 1727 8.127e-14
C404 1415 1727 6.946e-14
C402 1417 1727 1.275e-13
C400 1419 1727 1.8635e-14
C398 1421 1727 2.871e-14
C397 1422 1727 2.005e-14
C395 1424 1727 2.632e-14
C394 1425 1727 1.2482e-13
C393 1426 1727 2.321e-14
C391 1428 1727 5.165e-14
C390 1429 1727 4.869e-14
C381 1438 1727 7.43e-15
C379 1440 1727 9.7e-15
C377 1442 1727 1.0884e-13
C366 1453 1727 6.781e-14
C358 1461 1727 7.76e-15
C354 1465 1727 8.58e-15
C352 1467 1727 4.11e-15
C351 1468 1727 4.449e-14
C344 1474 1727 4.843e-14
C343 1475 1727 2.871e-14
C342 1476 1727 2.632e-14
C341 1477 1727 2.005e-14
C339 1479 1727 4.869e-14
C338 1480 1727 2.321e-14
C334 1484 1727 5.165e-14
C333 1485 1727 1.3671e-13
C332 1486 1727 2.445e-14
C331 1487 1727 5.474e-14
C329 1489 1727 5.281e-14
C327 1491 1727 2.596e-14
C326 1492 1727 2.16e-14
C323 1495 1727 5.725e-14
C321 1497 1727 1.677e-14
C320 1498 1727 9.204e-14
C319 1499 1727 1.8635e-14
C318 1500 1727 9.208e-14
C317 1501 1727 5.563e-14
C316 1502 1727 9.036e-14
C315 1503 1727 1.8635e-14
C314 1504 1727 9.446e-14
C313 1505 1727 7.43e-15
C312 1506 1727 4.151e-14
C310 1508 1727 9.183e-14
C308 1510 1727 2.871e-14
C305 1513 1727 4.869e-14
C304 1514 1727 2.321e-14
C303 1515 1727 2.632e-14
C301 1517 1727 2.005e-14
C300 1518 1727 5.165e-14
C299 1519 1727 7.458e-14
C298 1520 1727 7.155e-14
C295 1523 1727 5.356e-14
C294 1524 1727 5.346e-14
C290 1528 1727 6.761e-14
C288 1530 1727 8.34e-14
C287 1531 1727 2.596e-14
C286 1532 1727 2.16e-14
C283 1535 1727 5.169e-14
C282 1536 1727 1.1292e-13
C281 1537 1727 4.11e-15
C280 1538 1727 5.552e-14
C279 1539 1727 2.299e-14
C276 1542 1727 2.871e-14
C275 1543 1727 4.4277e-13
C274 1544 1727 2.632e-14
C273 1545 1727 4.869e-14
C271 1547 1727 2.005e-14
C270 1548 1727 5.165e-14
C269 1549 1727 2.321e-14
C268 1550 1727 7.69e-14
C265 1552 1727 2.871e-14
C263 1554 1727 2.005e-14
C261 1556 1727 2.632e-14
C259 1558 1727 5.165e-14
C258 1559 1727 2.321e-14
C257 1560 1727 4.869e-14
C256 1561 1727 1.767e-14
C255 1562 1727 5.598e-14
C254 1563 1727 6.05e-15
C253 1564 1727 5.981e-14
C252 1565 1727 2.605e-14
C250 1567 1727 5.411e-14
C249 1568 1727 1.8635e-14
C248 1569 1727 3.7539e-13
C247 1570 1727 1.6428e-13
C243 1574 1727 1.8128e-13
C242 1575 1727 8.529e-14
C241 1576 1727 1.568e-14
C240 1577 1727 1.8635e-14
C239 1578 1727 1.4695e-13
C238 1579 1727 8.452e-14
C237 1580 1727 2.605e-14
C236 1581 1727 3.5204e-13
C235 1582 1727 1.3795e-13
C234 1583 1727 1.8635e-14
C232 1585 1727 2.4639e-13
C231 1586 1727 3.8326e-13
C230 1587 1727 5.511e-14
C227 1590 1727 8.17e-14
C225 1592 1727 1.8635e-14
C223 1594 1727 9.02e-14
C222 1595 1727 1.8635e-14
C221 1596 1727 6.851e-14
C220 1597 1727 6.05e-15
C219 1598 1727 4.312e-14
C218 1599 1727 1.8635e-14
C217 1600 1727 4.873e-14
C216 1601 1727 4.17731e-13
C215 1602 1727 1.6884e-13
C214 1603 1727 1.8635e-14
C212 1605 1727 1.1836e-13
C211 1606 1727 1.8635e-14
C210 1607 1727 9.835e-14
C203 1614 1727 9.7e-15
C202 1615 1727 7.43e-15
C191 1626 1727 6.05e-15
C190 1627 1727 6.05e-15
C187 1629 1727 2.005e-14
C186 1630 1727 2.871e-14
C183 1633 1727 2.321e-14
C181 1635 1727 2.632e-14
C177 1639 1727 5.165e-14
C176 1640 1727 4.869e-14
C175 1641 1727 9.523e-14
C172 1644 1727 1.932e-14
C170 1646 1727 1.3654e-13
C167 1649 1727 2.356e-14
C166 1650 1727 1.4394e-13
C165 1651 1727 1.568e-14
C162 1654 1727 1.4796e-13
C161 1655 1727 1.568e-14
C159 1657 1727 6.249e-14
C158 1658 1727 2.596e-14
C156 1660 1727 2.16e-14
C152 1664 1727 5.725e-14
C151 1665 1727 2.445e-14
C146 1670 1727 5.401e-14
C144 1672 1727 7.945e-14
C143 1673 1727 5.233e-14
C142 1674 1727 1.8635e-14
C140 1676 1727 4.11e-15
C139 1677 1727 1.8525e-13
C135 1681 1727 2.005e-14
C132 1684 1727 2.632e-14
C130 1686 1727 2.871e-14
C129 1687 1727 9.314e-14
C128 1688 1727 2.321e-14
C127 1689 1727 4.869e-14
C126 1690 1727 5.165e-14
C123 1693 1727 1.8635e-14
C121 1695 1727 5.203e-14
C120 1696 1727 9.965e-14
C119 1697 1727 2.455e-14
C115 1701 1727 4.791e-14
C112 1704 1727 1.8635e-14
C109 1707 1727 5.203e-14
C108 1708 1727 1.81064e-12
C107 1709 1727 2.3741e-13
C106 1710 1727 6.33059e-13
C105 1711 1727 2.455e-14
C103 1713 1727 4.11e-15
C102 1714 1727 4.11e-15
C101 1715 1727 1.0786e-13
C100 1716 1727 6.947e-14
C97 1719 1727 5.621e-14
C95 1721 1727 1.767e-14
C94 1722 1727 4.727e-14
C92 1724 1727 1.8635e-14
C90 1726 1727 5.617e-14
C89 1727 1727 2.01874e-11
C88 1728 1727 8.155e-14
C86 1730 1727 2.871e-14
C85 1731 1727 2.005e-14
C83 1733 1727 2.321e-14
C81 1735 1727 2.632e-14
C80 1736 1727 5.358e-14
C79 1737 1727 5.165e-14
C78 1738 1727 4.869e-14
C77 1739 1727 5.141e-14
C76 1740 1727 6.05e-15
C75 1741 1727 1.767e-14
C74 1742 1727 5.741e-14
C73 1743 1727 2.605e-14
C70 1746 1727 2.871e-14
C69 1747 1727 2.005e-14
C68 1748 1727 4.869e-14
C67 1749 1727 2.321e-14
C65 1751 1727 2.632e-14
C64 1752 1727 2.1201e-13
C63 1753 1727 5.165e-14
C62 1754 1727 2.596e-14
C61 1755 1727 2.16e-14
C60 1756 1727 9.7e-15
C59 1757 1727 5.11e-14
C58 1758 1727 1.34768e-12
C57 1759 1727 7.278e-14
C56 1760 1727 6.05e-15
C55 1761 1727 1.767e-14
C54 1762 1727 6.735e-14
C52 1764 1727 4.577e-14
C51 1765 1727 7.181e-14
C50 1766 1727 4.449e-14
C49 1767 1727 8.958e-14
C48 1768 1727 2.605e-14
C47 1769 1727 2.6263e-13
C46 1770 1727 5.001e-14
C45 1771 1727 8.77099e-13
C44 1772 1727 8.73769e-13
C41 1775 1727 2.455e-14
C40 1776 1727 4.5038e-13
C39 1777 1727 1.8635e-14
C38 1778 1727 1.2786e-13
C36 1780 1727 8.005e-14
C35 1781 1727 7.378e-14
C34 1782 1727 1.8635e-14
C33 1783 1727 4.3732e-13
C32 1784 1727 6.591e-14
C31 1785 1727 5.2711e-13
C30 1786 1727 6.3355e-13
C29 1787 1727 2.596e-14
C28 1788 1727 2.16e-14
C27 1789 1727 9.7e-15
C26 1790 1727 1.4762e-13
C25 1791 1727 9.347e-14
C24 1792 1727 2.9748e-13
C23 1793 1727 6.915e-14
C22 1794 1727 6.05e-15
C21 1795 1727 4.432e-14
C20 1796 1727 5.692e-14
C19 1797 1727 6.31e-14
C18 1798 1727 2.299e-14
C16 1800 1727 8.58e-15
C15 1801 1727 1.1278e-13
C14 1802 1727 4.449e-14
C12 1804 1727 2.871e-14
C11 1805 1727 2.005e-14
C9 1807 1727 2.632e-14
C8 1808 1727 7.0871e-13
C7 1809 1727 7.69e-14
C6 1810 1727 2.76613e-12
C4 1812 1727 2.321e-14
C3 1813 1727 4.869e-14
C2 1814 1727 2.11053e-11
C1 1815 1727 5.165e-14
.ends act5_cougar

