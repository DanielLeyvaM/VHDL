* Spice description of mul5b_cougar
* Spice driver version -1209024860
* Date ( dd/mm/yyyy hh:mm:ss ): 28/10/2020 at 15:56:22

* INTERF vdd vss x[0] x[1] x[2] x[3] x[4] y[0] y[1] y[2] y[3] y[4] z[0] z[1] 
* INTERF z[2] z[3] z[4] z[5] z[6] z[7] z[8] z[9] 


.subckt mul5b_cougar 2127 2044 2113 2108 2125 2122 2123 2055 2058 1849 1457 1541 1933 1735 1538 1194 1446 1243 1120 480 235 567 
* NET 18 = xr2_x1_3_sig
* NET 23 = a2_x2_25_sig
* NET 24 = nao22_x1_37_sig
* NET 27 = na3_x1_22_sig
* NET 31 = na2_x1_35_sig
* NET 34 = na2_x1_33_sig
* NET 36 = na3_x1_23_sig
* NET 41 = on12_x1_6_sig
* NET 42 = aux6
* NET 44 = na4_x1_7_sig
* NET 48 = nao22_x1_40_sig
* NET 49 = ao22_x2_31_sig
* NET 52 = a2_x2_28_sig
* NET 57 = mx2_x2_6_sig
* NET 61 = aux214
* NET 62 = a3_x2_11_sig
* NET 69 = aux213
* NET 71 = na3_x1_24_sig
* NET 74 = na3_x1_25_sig
* NET 77 = o3_x2_10_sig
* NET 107 = not_aux8
* NET 110 = aux4
* NET 113 = ao22_x2_30_sig
* NET 116 = inv_x2_36_sig
* NET 117 = nao22_x1_38_sig
* NET 119 = a2_x2_26_sig
* NET 122 = not_aux211
* NET 126 = aux217
* NET 128 = on12_x1_4_sig
* NET 129 = no2_x1_17_sig
* NET 130 = na3_x1_21_sig
* NET 131 = na3_x1_20_sig
* NET 134 = ao22_x2_29_sig
* NET 137 = inv_x2_35_sig
* NET 138 = oa22_x2_19_sig
* NET 141 = na2_x1_34_sig
* NET 143 = nao22_x1_36_sig
* NET 144 = o3_x2_9_sig
* NET 148 = na3_x1_26_sig
* NET 149 = inv_x2_34_sig
* NET 150 = aux101
* NET 152 = na2_x1_31_sig
* NET 154 = nao22_x1_39_sig
* NET 155 = aux212
* NET 162 = inv_x2_5_sig
* NET 167 = a2_x2_3_sig
* NET 168 = aux5
* NET 169 = nao22_x1_sig
* NET 173 = inv_x2_4_sig
* NET 179 = aux198
* NET 182 = na4_x1_6_sig
* NET 184 = noa22_x1_13_sig
* NET 186 = na2_x1_36_sig
* NET 195 = not_aux6
* NET 198 = not_aux195
* NET 199 = ao22_x2_26_sig
* NET 200 = inv_x2_31_sig
* NET 205 = aux180
* NET 206 = aux181
* NET 214 = not_aux197
* NET 217 = inv_x2_33_sig
* NET 220 = noa22_x1_12_sig
* NET 221 = a4_x2_3_sig
* NET 230 = aux184
* NET 235 = z[8]
* NET 266 = not_aux227
* NET 272 = not_aux3
* NET 273 = inv_x2_3_sig
* NET 279 = a3_x2_10_sig
* NET 280 = no4_x1_2_sig
* NET 281 = a2_x2_27_sig
* NET 286 = no4_x1_3_sig
* NET 287 = a2_x2_24_sig
* NET 290 = nao22_x1_35_sig
* NET 291 = o2_x2_18_sig
* NET 295 = o3_x2_8_sig
* NET 296 = na2_x1_28_sig
* NET 297 = na3_x1_17_sig
* NET 298 = na4_x1_4_sig
* NET 301 = oa22_x2_16_sig
* NET 304 = not_aux225
* NET 305 = a2_x2_29_sig
* NET 308 = aux98
* NET 310 = not_aux149
* NET 313 = an12_x1_9_sig
* NET 315 = nao22_x1_34_sig
* NET 316 = nao22_x1_33_sig
* NET 317 = na4_x1_5_sig
* NET 318 = na2_x1_30_sig
* NET 319 = o2_x2_16_sig
* NET 320 = na3_x1_18_sig
* NET 323 = no2_x1_15_sig
* NET 324 = na3_x1_19_sig
* NET 325 = o2_x2_17_sig
* NET 330 = oa22_x2_17_sig
* NET 334 = not_aux1
* NET 343 = na2_x1_29_sig
* NET 345 = no4_x1_sig
* NET 348 = oa2a22_x2_6_sig
* NET 355 = not_aux154
* NET 359 = no2_x1_18_sig
* NET 362 = not_aux210
* NET 363 = aux207
* NET 368 = inv_x2_32_sig
* NET 377 = oa2ao222_x2_sig
* NET 381 = inv_x2_2_sig
* NET 386 = not_aux194
* NET 389 = not_aux23
* NET 390 = not_aux222
* NET 396 = a2_x2_23_sig
* NET 399 = a3_x2_9_sig
* NET 410 = xr2_x1_4_sig
* NET 411 = aux216
* NET 416 = a2_x2_21_sig
* NET 423 = aux87
* NET 429 = aux210
* NET 433 = na3_x1_16_sig
* NET 434 = na3_x1_15_sig
* NET 438 = ao22_x2_28_sig
* NET 443 = na2_x1_5_sig
* NET 452 = xr2_x1_6_sig
* NET 453 = aux29
* NET 457 = aux47
* NET 461 = no2_x1_19_sig
* NET 464 = no3_x1_4_sig
* NET 465 = aux61
* NET 468 = na2_x1_37_sig
* NET 469 = on12_x1_5_sig
* NET 474 = aux223
* NET 476 = nao22_x1_24_sig
* NET 477 = ao2o22_x2_sig
* NET 479 = oa22_x2_14_sig
* NET 480 = z[7]
* NET 488 = oa2a22_x2_5_sig
* NET 491 = o3_x2_7_sig
* NET 494 = o3_x2_6_sig
* NET 495 = no3_x1_2_sig
* NET 497 = oa22_x2_12_sig
* NET 498 = no2_x1_14_sig
* NET 501 = ao22_x2_27_sig
* NET 502 = na2_x1_26_sig
* NET 503 = na3_x1_14_sig
* NET 507 = no3_x1_3_sig
* NET 511 = noa2ao222_x1_sig
* NET 512 = na3_x1_13_sig
* NET 515 = an12_x1_8_sig
* NET 516 = no2_x1_13_sig
* NET 518 = na2_x1_27_sig
* NET 519 = not_aux208
* NET 522 = o2_x2_15_sig
* NET 524 = noa22_x1_11_sig
* NET 525 = nao22_x1_32_sig
* NET 527 = aux204
* NET 529 = a3_x2_8_sig
* NET 560 = a3_x2_12_sig
* NET 563 = o4_x2_sig
* NET 566 = noa22_x1_14_sig
* NET 567 = z[9]
* NET 574 = noa2ao222_x1_2_sig
* NET 576 = aux23
* NET 578 = oa22_x2_18_sig
* NET 579 = nao22_x1_42_sig
* NET 580 = ao22_x2_32_sig
* NET 583 = not_aux196
* NET 588 = not_aux209
* NET 589 = no3_x1_5_sig
* NET 590 = no2_x1_20_sig
* NET 596 = oa22_x2_15_sig
* NET 598 = aux177
* NET 600 = na3_x1_8_sig
* NET 602 = a4_x2_sig
* NET 612 = aux202
* NET 618 = aux172
* NET 620 = not_aux224
* NET 621 = na4_x1_3_sig
* NET 623 = not_aux172
* NET 628 = oa22_x2_13_sig
* NET 634 = noa22_x1_7_sig
* NET 638 = o2_x2_8_sig
* NET 642 = na2_x1_10_sig
* NET 649 = aux88
* NET 650 = aux156
* NET 651 = nao22_x1_29_sig
* NET 656 = noa22_x1_9_sig
* NET 659 = na2_x1_24_sig
* NET 663 = not_aux203
* NET 664 = xr2_x1_2_sig
* NET 667 = aux26
* NET 668 = ao2o22_x2_2_sig
* NET 674 = o2_x2_19_sig
* NET 677 = oa22_x2_20_sig
* NET 681 = not_aux200
* NET 683 = not_aux199
* NET 684 = o2_x2_11_sig
* NET 686 = na2_x1_21_sig
* NET 689 = noa22_x1_8_sig
* NET 690 = nao22_x1_26_sig
* NET 691 = na3_x1_10_sig
* NET 692 = oa2a22_x2_3_sig
* NET 693 = na4_x1_2_sig
* NET 697 = a2_x2_19_sig
* NET 698 = mbk_buf_aux98
* NET 701 = o2_x2_10_sig
* NET 702 = na3_x1_9_sig
* NET 705 = na2_x1_20_sig
* NET 708 = o2_x2_7_sig
* NET 709 = na3_x1_3_sig
* NET 710 = o3_x2_5_sig
* NET 715 = aux102
* NET 716 = not_aux102
* NET 717 = a4_x2_2_sig
* NET 719 = na2_x1_23_sig
* NET 720 = not_aux95
* NET 750 = not_aux26
* NET 751 = a2_x2_30_sig
* NET 752 = nao22_x1_41_sig
* NET 754 = inv_x2_37_sig
* NET 755 = na2_x1_6_sig
* NET 756 = not_aux48
* NET 759 = no2_x1_16_sig
* NET 761 = na2_x1_32_sig
* NET 766 = not_aux47
* NET 770 = a3_x2_6_sig
* NET 771 = aux221
* NET 773 = aux90
* NET 780 = aux179
* NET 782 = not_aux226
* NET 785 = oa2a2a2a24_x2_sig
* NET 787 = nao22_x1_27_sig
* NET 788 = nao22_x1_28_sig
* NET 794 = on12_x1_2_sig
* NET 799 = nao22_x1_25_sig
* NET 802 = not_aux201
* NET 805 = nao2o22_x1_2_sig
* NET 806 = a3_x2_5_sig
* NET 807 = a3_x2_4_sig
* NET 814 = na3_x1_4_sig
* NET 818 = na2_x1_11_sig
* NET 820 = not_aux193
* NET 824 = o2_x2_2_sig
* NET 830 = o2_x2_3_sig
* NET 834 = na2_x1_15_sig
* NET 835 = not_aux157
* NET 843 = not_aux13
* NET 846 = na3_x1_6_sig
* NET 847 = nao22_x1_21_sig
* NET 848 = oa22_x2_11_sig
* NET 849 = o2_x2_9_sig
* NET 850 = na3_x1_5_sig
* NET 854 = na3_x1_12_sig
* NET 856 = not_aux156
* NET 858 = na2_x1_18_sig
* NET 859 = not_aux99
* NET 862 = na2_x1_12_sig
* NET 870 = o3_x2_4_sig
* NET 871 = not_aux25
* NET 874 = an12_x1_10_sig
* NET 879 = nao22_x1_43_sig
* NET 880 = no2_x1_21_sig
* NET 885 = no2_x1_11_sig
* NET 889 = aux91
* NET 893 = oa2a22_x2_4_sig
* NET 897 = o2_x2_12_sig
* NET 901 = no3_x1_sig
* NET 906 = not_aux88
* NET 911 = not_aux71
* NET 914 = mx2_x2_5_sig
* NET 918 = nao22_x1_19_sig
* NET 926 = aux71
* NET 935 = nxr2_x1_2_sig
* NET 939 = not_aux0
* NET 940 = aux0
* NET 947 = aux182
* NET 951 = aux84
* NET 956 = xr2_x1_sig
* NET 961 = inv_x2_20_sig
* NET 962 = a2_x2_14_sig
* NET 970 = a3_x2_3_sig
* NET 971 = a2_x2_22_sig
* NET 974 = na3_x1_11_sig
* NET 975 = oa2a22_x2_2_sig
* NET 979 = na4_x1_sig
* NET 984 = not_aux91
* NET 987 = a2_x2_15_sig
* NET 989 = not_aux72
* NET 993 = not_aux173
* NET 996 = o2_x2_13_sig
* NET 997 = not_aux34
* NET 1004 = aux135
* NET 1005 = not_aux136
* NET 1006 = aux89
* NET 1009 = oa2a22_x2_sig
* NET 1010 = mx3_x2_18_sig
* NET 1018 = not_aux98
* NET 1068 = oa22_x2_2_sig
* NET 1069 = xr2_x1_5_sig
* NET 1078 = aux13
* NET 1081 = not_aux14
* NET 1082 = nao22_x1_6_sig
* NET 1094 = inv_x2_15_sig
* NET 1096 = not_aux86
* NET 1099 = aux49
* NET 1107 = on12_x1_sig
* NET 1113 = na2_x1_22_sig
* NET 1118 = o2_x2_6_sig
* NET 1119 = not_aux74
* NET 1120 = z[6]
* NET 1128 = mx3_x2_21_sig
* NET 1138 = aux174
* NET 1142 = not_aux100
* NET 1143 = a2_x2_10_sig
* NET 1145 = no2_x1_9_sig
* NET 1150 = na2_x1_8_sig
* NET 1152 = a3_x2_2_sig
* NET 1153 = ao22_x2_24_sig
* NET 1162 = nao22_x1_15_sig
* NET 1164 = not_aux31
* NET 1168 = not_aux170
* NET 1170 = oa22_x2_5_sig
* NET 1175 = no2_x1_10_sig
* NET 1177 = aux175
* NET 1179 = oa22_x2_6_sig
* NET 1183 = aux131
* NET 1184 = a2_x2_2_sig
* NET 1187 = inv_x2_26_sig
* NET 1189 = not_aux92
* NET 1190 = aux128
* NET 1194 = z[3]
* NET 1197 = mx3_x2_sig
* NET 1198 = mx3_x2_2_sig
* NET 1204 = aux219
* NET 1205 = inv_x2_10_sig
* NET 1209 = na2_x1_4_sig
* NET 1211 = not_aux28
* NET 1213 = na2_x1_3_sig
* NET 1214 = noa22_x1_4_sig
* NET 1221 = a2_x2_9_sig
* NET 1222 = ao22_x2_20_sig
* NET 1225 = no2_x1_6_sig
* NET 1226 = inv_x2_16_sig
* NET 1228 = na2_x1_7_sig
* NET 1233 = mx3_x2_8_sig
* NET 1235 = mx2_x2_3_sig
* NET 1236 = oa2ao222_x2_3_sig
* NET 1243 = z[5]
* NET 1246 = mx3_x2_7_sig
* NET 1252 = mx3_x2_16_sig
* NET 1254 = mx3_x2_17_sig
* NET 1261 = mx3_x2_14_sig
* NET 1263 = oa3ao322_x2_sig
* NET 1270 = nao22_x1_14_sig
* NET 1273 = aux93
* NET 1275 = ao22_x2_sig
* NET 1276 = not_aux137
* NET 1279 = na2_x1_2_sig
* NET 1280 = aux187
* NET 1281 = no2_x1_sig
* NET 1282 = not_aux220
* NET 1284 = nao2o22_x1_sig
* NET 1287 = inv_x2_19_sig
* NET 1288 = nao22_x1_10_sig
* NET 1290 = not_aux168
* NET 1291 = inv_x2_17_sig
* NET 1293 = not_aux101
* NET 1294 = na2_x1_sig
* NET 1339 = mx3_x2_3_sig
* NET 1346 = aux27
* NET 1349 = oa22_x2_3_sig
* NET 1350 = oa2ao222_x2_2_sig
* NET 1351 = inv_x2_6_sig
* NET 1355 = inv_x2_9_sig
* NET 1358 = oa22_x2_4_sig
* NET 1359 = aux18
* NET 1360 = inv_x2_7_sig
* NET 1363 = a2_x2_4_sig
* NET 1365 = aux16
* NET 1373 = not_aux22
* NET 1378 = mx3_x2_9_sig
* NET 1384 = nao22_x1_8_sig
* NET 1391 = not_aux144
* NET 1393 = nao22_x1_18_sig
* NET 1394 = mx3_x2_11_sig
* NET 1395 = oa22_x2_7_sig
* NET 1398 = nao22_x1_11_sig
* NET 1401 = na2_x1_9_sig
* NET 1406 = oa22_x2_10_sig
* NET 1407 = inv_x2_25_sig
* NET 1417 = na2_x1_17_sig
* NET 1419 = not_aux87
* NET 1420 = mx3_x2_10_sig
* NET 1424 = oa2ao222_x2_4_sig
* NET 1428 = not_aux134
* NET 1429 = inv_x2_18_sig
* NET 1431 = not_aux160
* NET 1434 = aux150
* NET 1435 = nmx2_x1_sig
* NET 1439 = aux126
* NET 1440 = mx2_x2_4_sig
* NET 1441 = na2_x1_14_sig
* NET 1446 = z[4]
* NET 1453 = ao22_x2_9_sig
* NET 1456 = ao22_x2_8_sig
* NET 1457 = y[3]
* NET 1460 = ao22_x2_19_sig
* NET 1463 = ao22_x2_21_sig
* NET 1464 = not_aux2
* NET 1469 = noa22_x1_5_sig
* NET 1470 = not_aux15
* NET 1473 = aux145
* NET 1474 = inv_x2_23_sig
* NET 1477 = a2_x2_13_sig
* NET 1479 = oa22_x2_9_sig
* NET 1487 = mx3_x2_12_sig
* NET 1488 = mx3_x2_13_sig
* NET 1492 = oa2ao222_x2_5_sig
* NET 1499 = nao22_x1_12_sig
* NET 1504 = nao22_x1_20_sig
* NET 1505 = mx3_x2_19_sig
* NET 1508 = mx3_x2_20_sig
* NET 1515 = na2_x1_16_sig
* NET 1517 = nao22_x1_31_sig
* NET 1522 = aux147
* NET 1524 = an12_x1_6_sig
* NET 1527 = not_aux164
* NET 1529 = o2_x2_sig
* NET 1532 = o2_x2_14_sig
* NET 1533 = not_aux126
* NET 1537 = inv_x2_sig
* NET 1538 = z[2]
* NET 1539 = nao22_x1_3_sig
* NET 1540 = nao22_x1_2_sig
* NET 1541 = y[4]
* NET 1542 = ao22_x2_7_sig
* NET 1544 = not_y[4]
* NET 1546 = ao22_x2_18_sig
* NET 1553 = not_aux17
* NET 1567 = not_aux161
* NET 1569 = inv_x2_29_sig
* NET 1570 = not_aux167
* NET 1577 = not_aux206
* NET 1579 = inv_x2_27_sig
* NET 1581 = not_aux179
* NET 1596 = no2_x1_2_sig
* NET 1599 = ao22_x2_15_sig
* NET 1600 = ao22_x2_13_sig
* NET 1603 = ao22_x2_14_sig
* NET 1607 = no2_x1_3_sig
* NET 1608 = inv_x2_8_sig
* NET 1609 = not_aux218
* NET 1610 = not_aux20
* NET 1616 = inv_x2_13_sig
* NET 1620 = mx3_x2_6_sig
* NET 1624 = mx2_x2_sig
* NET 1628 = ao22_x2_16_sig
* NET 1629 = not_aux76
* NET 1632 = not_aux40
* NET 1634 = noa22_x1_3_sig
* NET 1637 = oa2ao222_x2_7_sig
* NET 1638 = inv_x2_24_sig
* NET 1642 = a2_x2_17_sig
* NET 1645 = noa22_x1_6_sig
* NET 1648 = ao22_x2_25_sig
* NET 1651 = oa2ao222_x2_9_sig
* NET 1653 = not_aux143
* NET 1654 = not_aux176
* NET 1656 = aux186
* NET 1657 = nao22_x1_13_sig
* NET 1658 = not_aux39
* NET 1661 = nao22_x1_17_sig
* NET 1662 = mx3_x2_15_sig
* NET 1665 = nao22_x1_16_sig
* NET 1673 = not_aux184
* NET 1674 = no2_x1_12_sig
* NET 1676 = nao22_x1_30_sig
* NET 1677 = oa2ao222_x2_8_sig
* NET 1678 = inv_x2_28_sig
* NET 1682 = not_aux190
* NET 1683 = na2_x1_13_sig
* NET 1684 = aux192
* NET 1685 = a2_x2_18_sig
* NET 1689 = an12_x1_5_sig
* NET 1714 = aux118
* NET 1721 = oa2ao222_x2_6_sig
* NET 1735 = z[1]
* NET 1739 = ao22_x2_2_sig
* NET 1742 = ao22_x2_5_sig
* NET 1745 = a3_x2_sig
* NET 1747 = aux30
* NET 1749 = o3_x2_3_sig
* NET 1753 = not_y[0]
* NET 1754 = ao22_x2_23_sig
* NET 1755 = o3_x2_2_sig
* NET 1757 = not_y[3]
* NET 1759 = mx3_x2_5_sig
* NET 1762 = mx3_x2_4_sig
* NET 1763 = nao22_x1_5_sig
* NET 1764 = not_y[2]
* NET 1769 = nmx3_x1_sig
* NET 1772 = inv_x2_12_sig
* NET 1776 = inv_x2_11_sig
* NET 1783 = o3_x2_sig
* NET 1784 = nao22_x1_4_sig
* NET 1789 = not_aux83
* NET 1791 = inv_x2_22_sig
* NET 1792 = not_aux9
* NET 1793 = oa22_x2_8_sig
* NET 1795 = not_aux68
* NET 1796 = not_aux70
* NET 1799 = na3_x1_2_sig
* NET 1802 = a2_x2_16_sig
* NET 1807 = not_aux104
* NET 1809 = not_aux146
* NET 1812 = a2_x2_20_sig
* NET 1816 = a3_x2_7_sig
* NET 1817 = nao22_x1_22_sig
* NET 1820 = na2_x1_19_sig
* NET 1821 = on12_x1_3_sig
* NET 1822 = na3_x1_7_sig
* NET 1827 = not_aux90
* NET 1831 = not_aux191
* NET 1839 = ao22_x2_3_sig
* NET 1842 = not_aux56
* NET 1843 = noa22_x1_sig
* NET 1848 = ao22_x2_11_sig
* NET 1849 = y[2]
* NET 1852 = not_aux55
* NET 1853 = noa22_x1_2_sig
* NET 1855 = na3_x1_sig
* NET 1858 = ao22_x2_22_sig
* NET 1860 = no2_x1_7_sig
* NET 1864 = not_aux46
* NET 1866 = no2_x1_8_sig
* NET 1867 = mx2_x2_2_sig
* NET 1872 = inv_x2_14_sig
* NET 1873 = not_aux78
* NET 1877 = not_aux165
* NET 1878 = aux94
* NET 1880 = inv_x2_30_sig
* NET 1881 = nao22_x1_23_sig
* NET 1883 = inv_x2_21_sig
* NET 1884 = not_y[1]
* NET 1885 = not_aux117
* NET 1886 = oa22_x2_sig
* NET 1891 = nao22_x1_7_sig
* NET 1893 = not_aux105
* NET 1895 = a2_x2_12_sig
* NET 1896 = nao22_x1_9_sig
* NET 1898 = not_x[3]
* NET 1899 = not_x[4]
* NET 1900 = not_aux103
* NET 1901 = aux183
* NET 1902 = na2_x1_25_sig
* NET 1903 = noa22_x1_10_sig
* NET 1907 = aux103
* NET 1933 = z[0]
* NET 1935 = aux50
* NET 1940 = an12_x1_2_sig
* NET 1941 = ao22_x2_6_sig
* NET 1947 = a2_x2_6_sig
* NET 1948 = a2_x2_8_sig
* NET 1949 = ao22_x2_12_sig
* NET 1954 = an12_x1_4_sig
* NET 1956 = aux215
* NET 1962 = aux20
* NET 1966 = aux53
* NET 1972 = ao22_x2_17_sig
* NET 1973 = no2_x1_5_sig
* NET 1976 = no2_x1_4_sig
* NET 1977 = not_aux38
* NET 1981 = not_aux12
* NET 1984 = an12_x1_7_sig
* NET 1988 = aux81
* NET 1994 = not_aux77
* NET 1995 = not_aux79
* NET 2001 = nxr2_x1_sig
* NET 2010 = aux10
* NET 2011 = a2_x2_11_sig
* NET 2014 = not_aux125
* NET 2015 = a2_x2_sig
* NET 2019 = aux62
* NET 2022 = not_aux63
* NET 2028 = not_aux115
* NET 2029 = not_aux110
* NET 2030 = o2_x2_5_sig
* NET 2036 = not_aux121
* NET 2039 = not_aux124
* NET 2041 = not_aux109
* NET 2043 = o2_x2_4_sig
* NET 2044 = vss
* NET 2045 = ao22_x2_4_sig
* NET 2048 = an12_x1_sig
* NET 2049 = a2_x2_5_sig
* NET 2055 = y[0]
* NET 2056 = ao22_x2_10_sig
* NET 2058 = y[1]
* NET 2059 = an12_x1_3_sig
* NET 2062 = a2_x2_7_sig
* NET 2063 = aux60
* NET 2066 = aux19
* NET 2069 = not_aux45
* NET 2070 = aux59
* NET 2074 = not_aux44
* NET 2075 = not_aux43
* NET 2079 = not_aux37
* NET 2083 = not_aux35
* NET 2087 = aux34
* NET 2088 = mbk_buf_aux34
* NET 2092 = not_aux33
* NET 2093 = not_aux64
* NET 2095 = aux66
* NET 2096 = not_aux66
* NET 2098 = not_aux32
* NET 2101 = mbk_buf_aux31
* NET 2102 = aux31
* NET 2104 = not_aux106
* NET 2105 = not_x[1]
* NET 2108 = x[1]
* NET 2109 = not_aux171
* NET 2111 = not_aux67
* NET 2113 = x[0]
* NET 2115 = not_x[0]
* NET 2119 = not_aux112
* NET 2120 = aux111
* NET 2121 = not_aux111
* NET 2122 = x[3]
* NET 2123 = x[4]
* NET 2125 = x[2]
* NET 2126 = not_x[2]
* NET 2127 = vdd
Mtr_04128 2120 2124 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04127 2127 2122 2124 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04126 2124 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04125 2126 2125 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04124 2127 2125 2126 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04123 2127 2125 2126 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04122 2126 2125 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04121 2127 2116 2118 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04120 2118 2117 2119 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04119 2118 2120 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04118 2119 2125 2118 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04117 2127 2120 2117 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04116 2116 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04115 2121 2120 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04114 2101 2103 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04113 2127 2102 2103 2127 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_04112 2106 2105 2107 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04111 2127 2111 2106 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04110 2104 2107 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04109 2109 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04108 2127 2111 2109 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04107 2127 2110 2112 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04106 2112 2114 2111 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04105 2112 2125 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04104 2111 2123 2112 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04103 2127 2125 2114 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04102 2110 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04101 2127 2113 2094 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04100 2095 2093 2094 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04099 2094 2092 2095 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04098 2097 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04097 2127 2102 2100 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04096 2098 2097 2099 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04095 2099 2102 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04094 2099 2100 2098 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04093 2127 2123 2099 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04092 2096 2095 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04091 2115 2113 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04090 2102 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04089 2127 2126 2102 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04088 2086 2126 2087 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04087 2127 2122 2086 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04086 2088 2089 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04085 2127 2087 2089 2127 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_04084 2077 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04083 2076 2098 2078 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04082 2127 2105 2076 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04081 2078 2083 2077 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04080 2075 2078 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04079 2127 2080 2079 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04078 2080 2092 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04077 2127 2105 2081 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04076 2081 2083 2080 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04075 2127 2082 2085 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04074 2085 2084 2083 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04073 2085 2087 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04072 2083 2123 2085 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04071 2127 2087 2084 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04070 2082 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04069 2091 2098 2090 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04068 2127 2108 2091 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04067 2092 2090 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04066 2127 2065 2068 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04065 2068 2067 2069 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04064 2068 2066 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04063 2069 2123 2068 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04062 2127 2066 2067 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04061 2065 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04060 2063 2064 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04059 2127 2069 2064 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04058 2064 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04057 2070 2071 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04056 2127 2075 2071 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04055 2071 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04054 2073 2115 2072 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04053 2127 2075 2073 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04052 2074 2072 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04051 2049 2054 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04050 2127 2063 2054 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04049 2054 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04048 2046 2070 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04047 2127 2046 2047 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04046 2047 2058 2048 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04045 2052 2063 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04044 2127 2052 2053 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04043 2053 2058 2059 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04042 2127 2057 2056 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04041 2057 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04040 2127 2059 2061 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04039 2061 2062 2057 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04038 2062 2060 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04037 2127 2070 2060 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04036 2060 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04035 2127 2050 2045 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04034 2050 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04033 2127 2048 2051 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04032 2051 2049 2050 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04031 1932 2105 2042 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04030 2127 2041 1932 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04029 2043 2042 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04028 1930 2119 2035 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04027 2127 2108 1930 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04026 2036 2035 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04025 2127 2037 2039 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04024 1931 2115 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04023 1931 2043 2037 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04022 2037 2036 1931 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04021 1929 2105 2033 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04020 2127 2119 1929 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_04019 2030 2033 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04018 2127 2026 2028 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04017 1928 2115 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04016 1928 2030 2026 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04015 2026 2029 1928 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04014 2127 2017 2014 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04013 2017 2039 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04012 2127 2015 1926 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04011 1926 2113 2017 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04010 2011 2013 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04009 2127 2010 2013 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04008 2013 2109 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04007 2127 2020 1927 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04006 1927 2027 2022 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04005 1927 2019 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04004 2022 2123 1927 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04003 2127 2019 2027 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04002 2020 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_04001 2015 2008 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_04000 2127 2010 2008 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03999 2008 2104 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03998 1923 2105 1997 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03997 2127 2022 1923 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03996 2093 1997 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03995 2127 2113 1921 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03994 1988 1995 1921 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03993 1921 2092 1988 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03992 1995 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03991 2127 2022 1995 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03990 2127 2000 1924 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03989 1924 2002 2001 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03988 1924 2010 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03987 2001 2122 1924 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03986 2127 2010 2002 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03985 2000 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03984 1925 2126 2006 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03983 2127 2108 1925 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03982 2010 2006 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03981 2127 1990 1922 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03980 1922 1992 1994 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03979 1922 2123 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03978 1994 2108 1922 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03977 2127 2123 1992 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03976 1990 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03975 2127 1974 1972 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03974 1974 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03973 2127 1973 1917 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03972 1917 1976 1974 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03971 2127 2001 1981 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03970 1981 1980 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03969 2127 2113 1980 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03968 1919 2115 1978 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03967 2127 2079 1919 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03966 1977 1978 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03965 1985 2074 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03964 2127 1985 1920 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03963 1920 1988 1984 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03962 1918 2074 1976 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03961 2127 2058 1918 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03960 1947 1946 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03959 2127 1966 1946 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03958 1946 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03957 1963 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03956 2127 2122 1967 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03955 2066 1963 1916 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03954 1916 2122 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03953 1916 1967 2066 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03952 2127 2108 1916 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03951 1956 1958 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03950 2127 2113 1958 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03949 1958 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03948 1966 1970 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03947 2127 2079 1970 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03946 1970 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03945 1955 1966 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03944 2127 1955 1914 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03943 1914 2058 1954 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03942 1960 2066 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03941 2127 1960 1915 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03940 1915 2113 1962 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03939 1938 1935 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03938 2127 1938 1911 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03937 1911 2058 1940 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03936 1933 1934 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03935 2127 1956 1934 2127 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_03934 2127 1950 1949 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03933 1950 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03932 2127 1948 1913 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03931 1913 1954 1950 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03930 1948 1936 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03929 2127 1935 1936 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03928 1936 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03927 2127 1942 1941 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03926 1942 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03925 2127 1940 1912 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03924 1912 1947 1942 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03923 2127 1908 1910 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03922 1910 1909 2041 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03921 1910 1907 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03920 2041 2125 1910 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03919 2127 1907 1909 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03918 1908 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03917 1900 1907 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03916 2127 2115 1905 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03915 1903 1902 1905 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03914 1905 2029 1903 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03913 1902 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03912 2127 1901 1902 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03911 1904 2041 1906 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03910 2127 2108 1904 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03909 2029 1906 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03908 2127 2028 1891 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03907 1892 2113 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03906 1891 2011 1892 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03905 2127 1887 1885 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03904 1888 1884 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03903 1888 1886 1887 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03902 1887 2028 1888 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03901 2127 2039 1896 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03900 1897 2113 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03899 1896 1895 1897 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03898 1907 1899 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03897 2127 1898 1907 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03896 2127 1889 1886 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03895 1890 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03894 1890 2104 1889 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03893 1889 1893 1890 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03892 1895 1894 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03891 2127 2109 1894 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03890 1894 1893 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03889 1899 2123 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03888 2127 2123 1899 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03887 2127 2123 1899 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03886 1899 2123 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03885 1883 1885 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03884 1876 2115 1879 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03883 2127 1994 1876 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03882 1877 1879 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03881 1880 1878 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03880 2127 1885 1881 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03879 1882 2058 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03878 1881 1880 1882 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03877 1865 1884 1973 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03876 2127 1864 1865 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03875 1878 2096 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03874 2127 1977 1878 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03873 2127 1871 1867 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03872 1870 1988 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03871 1868 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03870 1869 2058 1871 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03869 1871 1868 1870 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03868 2127 1872 1869 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03867 1872 1873 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03866 1875 1994 1874 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03865 2127 2113 1875 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03864 1873 1874 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03863 1862 1884 1866 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03862 2127 2074 1862 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03861 1859 1864 1860 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03860 2127 2058 1859 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03859 1856 2115 1857 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03858 2127 2069 1856 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03857 1864 1857 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03856 2127 2058 1855 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03855 1855 1898 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03854 1855 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03853 2127 1863 1858 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03852 1863 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03851 2127 1866 1861 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03850 1861 1860 1863 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03849 2127 1850 1848 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03848 1850 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03847 2127 1949 1851 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03846 1851 1853 1850 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03845 2127 2055 1854 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03844 1853 1855 1854 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03843 1854 1852 1853 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03842 2127 2055 1844 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03841 1843 1852 1844 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03840 1844 1842 1843 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03839 1935 1838 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03838 2127 1899 1838 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03837 1838 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03836 2127 1841 1839 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03835 1841 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03834 2127 2045 1840 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03833 1840 1843 1841 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03832 2127 2125 1845 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03831 1845 2058 1846 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03830 1846 2115 1847 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03829 1852 1847 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03828 2127 1820 1822 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03827 1822 1821 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03826 1822 2115 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03825 2127 2105 1821 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03824 1821 1825 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03823 2127 1901 1825 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03822 2127 1827 1732 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03821 1901 2126 1732 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03820 1732 2121 1901 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03819 1733 2126 1830 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03818 2127 2121 1733 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03817 1831 1830 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03816 1832 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03815 2127 2125 1833 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03814 2019 1832 1734 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03813 1734 2125 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03812 1734 1833 2019 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03811 2127 2122 1734 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03810 2127 1822 1814 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03809 1816 1814 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03808 2127 1884 1814 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03807 1814 1817 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03806 1812 1808 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03805 2127 1809 1808 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03804 1808 1807 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03803 1726 1807 1803 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03802 2127 2108 1726 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03801 1893 1803 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03800 1727 1900 1805 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03799 2127 2125 1727 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03798 1807 1805 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03797 2127 2104 1817 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03796 1728 2108 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03795 1817 1812 1728 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03794 1721 1797 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03793 1723 1883 1722 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03792 1723 1753 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03791 2127 1793 1723 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03790 1722 1802 1797 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03789 1797 2055 1723 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03788 1802 1800 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03787 2127 1884 1800 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03786 1800 1799 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03785 2127 1794 1796 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03784 1719 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03783 1719 2093 1794 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03782 1794 1795 1719 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03781 2127 1790 1793 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03780 1717 1791 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03779 1717 1878 1790 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03778 1790 2058 1717 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03777 2127 1788 1789 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03776 1715 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03775 1715 1995 1788 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03774 1788 1795 1715 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03773 1707 1775 1780 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03772 2127 1773 1708 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03771 1706 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03770 1780 1784 1706 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03769 1708 1772 1707 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03768 1709 1776 1708 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03767 1780 1884 1709 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03766 1762 1780 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03765 1775 1884 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03764 2127 2055 1773 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03763 1714 1796 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03762 2127 2074 1714 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03761 2127 1783 1784 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03760 1710 1981 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03759 1784 1884 1710 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03758 2127 2113 1712 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03757 1712 2058 1711 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03756 1711 2126 1786 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03755 1783 1786 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03754 1791 1792 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03753 1772 1796 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03752 1702 1765 1769 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03751 2127 1758 1703 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03750 1701 1757 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03749 1769 1759 1701 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03748 1703 1763 1702 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03747 1704 1762 1703 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03746 1769 1764 1704 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03745 1765 1764 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03744 2127 1757 1758 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03743 2127 1755 1763 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03742 1699 1753 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03741 1763 1754 1699 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03740 2127 2113 1695 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03739 1695 2058 1696 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03738 1696 1899 1746 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03737 1749 1746 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03736 1705 1898 1771 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03735 2127 2058 1705 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03734 1792 1771 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03733 2127 1750 1754 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03732 1750 1749 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03731 2127 2096 1698 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03730 1698 1884 1750 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03729 2127 1741 1742 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03728 1741 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03727 2127 1941 1692 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03726 1692 1745 1741 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03725 1747 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03724 2127 2058 1747 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03723 2127 1753 1744 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03722 1745 1744 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03721 2127 1747 1744 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03720 1744 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03719 1736 1753 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03718 2127 1736 1688 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03717 1688 1747 1689 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03716 2127 1738 1739 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03715 1738 1757 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03714 2127 1742 1690 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03713 1690 1839 1738 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03712 1685 1686 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03711 2127 1684 1686 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03710 1686 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03709 1683 2036 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03708 2127 1682 1683 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03707 2127 2058 1676 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03706 1675 1674 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03705 1676 1903 1675 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03704 1820 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03703 2127 1673 1820 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03702 1677 1679 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03701 1681 1678 1680 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03700 1681 2115 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03699 2127 1683 1681 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03698 1680 1685 1679 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03697 1679 2113 1681 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03696 1678 1795 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03695 1668 1666 1667 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03694 2127 1663 1669 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03693 1664 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03692 1667 1661 1664 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03691 1669 1677 1668 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03690 1670 1665 1669 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03689 1667 2058 1670 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03688 1662 1667 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03687 1666 2058 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03686 2127 2055 1663 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03685 1672 2111 1671 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03684 2127 2108 1672 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03683 1795 1671 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03682 2127 1658 1661 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03681 1660 2014 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03680 1661 1884 1660 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03679 1636 2126 1635 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03678 2127 2058 1636 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03677 1658 1635 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03676 2127 2115 1644 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03675 1645 1795 1644 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03674 1644 1654 1645 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03673 2127 1653 1657 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03672 1659 2058 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03671 1657 2014 1659 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03670 1651 1650 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03669 1652 1648 1649 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03668 1652 1753 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03667 2127 1881 1652 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03666 1649 1816 1650 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03665 1650 2055 1652 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03664 2127 2113 1655 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03663 1656 1654 1655 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03662 1655 1893 1656 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03661 2127 1647 1648 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03660 1647 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03659 2127 1645 1646 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03658 1646 1656 1647 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03657 2127 2055 1633 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03656 1634 1632 1633 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03655 1633 1658 1634 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03654 2127 1631 1628 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03653 1631 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03652 2127 1972 1630 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03651 1630 1634 1631 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03650 1638 1658 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03649 1776 1629 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03648 1637 1639 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03647 1640 1638 1641 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03646 1640 2055 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03645 2127 1657 1640 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03644 1641 1642 1639 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03643 1639 1753 1640 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03642 1642 1643 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03641 2127 1714 1643 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03640 1643 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03639 2127 1615 1624 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03638 1614 1962 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03637 1617 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03636 1618 2058 1615 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03635 1615 1617 1614 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03634 2127 1616 1618 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03633 2127 2113 1611 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03632 1611 1609 1613 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03631 1613 1898 1612 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03630 1755 1612 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03629 1604 1884 1607 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03628 2127 1977 1604 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03627 1622 1625 1621 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03626 2127 1619 1626 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03625 1623 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03624 1621 1620 1623 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03623 1626 1867 1622 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03622 1627 1624 1626 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03621 1621 2055 1627 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03620 1759 1621 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03619 1625 2055 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03618 2127 1764 1619 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03617 1608 1792 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03616 1610 1962 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03615 2127 1598 1599 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03614 1598 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03613 2127 1607 1597 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03612 1597 1596 1598 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03611 2127 1601 1603 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03610 1601 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03609 2127 1599 1602 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03608 1602 1689 1601 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03607 2127 1605 1600 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03606 1605 1757 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03605 2127 1628 1606 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03604 1606 1603 1605 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03603 1595 1899 1596 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03602 2127 2058 1595 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03601 1537 1684 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03600 1531 1831 1589 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03599 2127 2108 1531 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03598 1532 1589 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03597 1684 1831 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03596 2127 1533 1684 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03595 1530 1577 1674 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03594 2127 2113 1530 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03593 2127 1592 1577 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03592 1592 1682 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03591 2127 1537 1535 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03590 1535 2108 1592 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03589 1521 2109 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03588 2127 1521 1523 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03587 1523 1522 1524 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03586 2127 2096 1517 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03585 1516 1577 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03584 1517 2115 1516 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03583 2127 1579 1665 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03582 1519 1581 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03581 1665 2111 1519 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03580 2127 1585 1527 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03579 1525 1529 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03578 1525 1900 1585 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03577 1585 2126 1525 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03576 1528 2113 1586 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03575 2127 2108 1528 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03574 1529 1586 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03573 1515 1581 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03572 2127 1527 1515 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03571 2127 1572 1570 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03570 1502 1884 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03569 1502 1877 1572 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03568 1572 1527 1502 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03567 2127 1570 1499 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03566 1497 2058 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03565 1499 1567 1497 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03564 1410 1513 1511 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03563 2127 1507 1411 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03562 1405 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03561 1511 1504 1405 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03560 1411 1508 1410 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03559 1409 1515 1411 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03558 1511 1884 1409 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03557 1505 1511 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03556 1513 1884 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03555 2127 2055 1507 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03554 2127 1570 1504 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03553 1500 2058 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03552 1504 1569 1500 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03551 1569 1473 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03550 1380 1494 1496 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03549 2127 1490 1389 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03548 1381 1757 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03547 1496 1488 1381 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03546 1389 1721 1380 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03545 1390 1492 1389 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03544 1496 1849 1390 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03543 1487 1496 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03542 1494 1849 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03541 2127 1757 1490 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03540 1372 1484 1482 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03539 2127 1481 1376 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03538 1371 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03537 1482 1637 1371 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03536 1376 1479 1372 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03535 1377 1499 1376 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03534 1482 1753 1377 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03533 1488 1482 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03532 1484 1753 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03531 2127 1849 1481 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03530 1473 1864 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03529 2127 1629 1473 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03528 1477 1560 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03527 2127 1864 1560 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03526 1560 1873 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03525 2127 1561 1479 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03524 1475 1474 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03523 1475 1473 1561 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03522 1561 2058 1475 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03521 1471 1884 1555 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03520 2127 1470 1471 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03519 1632 1555 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03518 1616 1464 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03517 2127 2055 1467 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03516 1469 1632 1467 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03515 1467 1553 1469 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03514 2127 1551 1463 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03513 1551 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03512 2127 1858 1465 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03511 1465 1469 1551 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03510 2127 1550 1546 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03509 1550 1457 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03508 2127 1463 1461 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03507 1461 1460 1550 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03506 2127 1539 1446 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03505 1446 1540 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03504 1446 1769 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03503 2127 1545 1456 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03502 1545 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03501 2127 2056 1454 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03500 1454 1453 1545 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03499 2127 1541 1540 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03498 1449 1542 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03497 1540 1739 1449 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03496 2127 1548 1542 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03495 1548 1457 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03494 2127 1848 1458 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03493 1458 1456 1548 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03492 2127 1544 1539 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03491 1451 1546 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03490 1539 1600 1451 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03489 2127 1444 1440 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03488 1443 1441 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03487 1445 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03486 1442 2108 1444 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03485 1444 1445 1443 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03484 2127 2019 1442 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03483 1533 1439 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03482 2127 1433 1567 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03481 1433 1431 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03480 2127 1435 1432 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03479 1432 2113 1433 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03478 1435 1438 1436 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03477 1437 2108 1435 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03476 1436 1434 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03475 2127 1522 1437 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03474 1438 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03473 1441 1533 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03472 2127 1673 1441 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03471 1429 1428 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03470 1426 1422 1427 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03469 2127 1423 1430 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03468 1421 1884 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03467 1427 1896 1421 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03466 1430 1424 1426 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03465 1425 1429 1430 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03464 1427 2115 1425 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03463 1420 1427 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03462 1422 2115 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03461 2127 1884 1423 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03460 1416 1412 1415 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03459 2127 1413 1418 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03458 1408 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03457 1415 1406 1408 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03456 1418 1417 1416 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03455 1414 1900 1418 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03454 1415 2105 1414 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03453 1508 1415 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03452 1412 2105 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03451 2127 2113 1413 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03450 1417 1673 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03449 2127 1899 1417 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03448 1522 1809 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03447 2127 2101 1522 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03446 1809 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03445 2127 1419 1809 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03444 1388 1382 1386 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03443 2127 1383 1387 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03442 1379 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03441 1386 1394 1379 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03440 1387 1420 1388 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03439 1385 1384 1387 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03438 1386 2055 1385 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03437 1378 1386 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03436 1382 2055 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03435 2127 1849 1383 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03434 1407 1714 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03433 1400 1396 1402 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03432 2127 1397 1403 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03431 1399 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03430 1402 1398 1399 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03429 1403 1395 1400 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03428 1404 1401 1403 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03427 1402 2058 1404 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03426 1394 1402 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03425 1396 2058 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03424 2127 2055 1397 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03423 1401 1877 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03422 2127 1464 1401 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03421 2127 1391 1393 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03420 1392 1567 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03419 1393 1884 1392 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03418 2127 1373 1384 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03417 1374 1884 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03416 1384 1984 1374 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03415 1474 1391 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03414 1367 2105 1368 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03413 2127 2058 1367 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03412 1553 1368 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03411 2127 1553 1398 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03410 1369 1477 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03409 1398 1884 1369 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03408 2127 1365 1391 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03407 1391 1366 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03406 2127 2058 1366 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03405 2127 1361 1358 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03404 1362 1360 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03403 1362 1359 1361 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03402 1361 2058 1362 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03401 1363 1364 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03400 2127 1365 1364 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03399 1364 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03398 1365 1470 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03397 2127 1981 1365 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03396 1360 1553 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03395 1370 2105 1375 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03394 2127 2113 1370 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03393 1464 1375 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03392 1355 1609 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03391 2127 1347 1349 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03390 1348 1351 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03389 1348 1346 1347 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03388 1347 2058 1348 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03387 2127 1356 1373 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03386 1357 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03385 1357 1470 1356 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03384 1356 1610 1357 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03383 1344 1341 1343 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03382 2127 1338 1345 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03381 1340 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03380 1343 1350 1340 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03379 1345 1358 1344 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03378 1342 1349 1345 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03377 1343 1753 1342 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03376 1339 1343 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03375 1341 1753 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03374 2127 1849 1338 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03373 1350 1352 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03372 1354 1608 1353 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03371 1354 2125 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03370 2127 1355 1354 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03369 1353 1363 1352 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03368 1352 2055 1354 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03367 1351 1373 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03366 2127 1290 1288 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03365 1181 2105 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03364 1288 1434 1181 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03363 1291 1290 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03362 1163 1428 1281 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03361 2127 1884 1163 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03360 2127 1295 1682 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03359 1193 2105 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03358 1193 1294 1295 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03357 1295 1293 1193 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03356 1294 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03355 2127 1900 1294 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03354 1186 1419 1439 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03353 2127 2125 1186 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03352 1287 1431 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03351 2127 1285 1395 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03350 1176 1287 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03349 1176 1288 1285 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03348 1285 2115 1176 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03347 2127 1281 1653 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03346 1159 1275 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03345 1653 1279 1159 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03344 1284 1524 1171 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03343 1171 2113 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03342 1167 1900 1284 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03341 2127 1282 1167 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03340 1279 1276 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03339 2127 2115 1279 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03338 1579 1280 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03337 2127 1653 1270 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03336 1156 2058 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03335 1270 1407 1156 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03334 1149 1269 1267 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03333 2127 1264 1148 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03332 1141 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03331 1267 1662 1141 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03330 1148 1263 1149 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03329 1147 1270 1148 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03328 1267 2055 1147 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03327 1261 1267 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03326 1269 2055 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03325 2127 1849 1264 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03324 2127 1272 1275 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03323 1272 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03322 2127 1273 1157 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03321 1157 1827 1272 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03320 1136 1260 1259 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03319 2127 1255 1137 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03318 1132 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03317 1259 1505 1132 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03316 1137 1254 1136 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03315 1135 1393 1137 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03314 1259 2055 1135 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03313 1252 1259 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03312 1260 2055 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03311 2127 1764 1255 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03310 1124 1249 1247 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03309 2127 1245 1125 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03308 1117 1541 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03307 1247 1487 1117 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03306 1125 1378 1124 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03305 1123 1246 1125 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03304 1247 1757 1123 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03303 1243 1247 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03302 1249 1757 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03301 2127 1541 1245 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03300 1228 1789 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03299 2127 1977 1228 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03298 2127 1231 1235 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03297 1104 1228 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03296 1229 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03295 1103 2058 1231 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03294 1231 1229 1104 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03293 2127 1359 1103 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03292 1226 1789 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03291 1115 1239 1241 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03290 2127 1237 1116 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03289 1112 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03288 1241 1233 1112 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03287 1116 1236 1115 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03286 1114 1235 1116 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03285 1241 2055 1114 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03284 1246 1241 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03283 1239 2055 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03282 2127 1764 1237 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03281 1098 1977 1225 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03280 2127 2058 1098 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03279 2127 1223 1222 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03278 1223 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03277 2127 1221 1095 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03276 1095 1225 1223 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03275 2127 1217 1092 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03274 1092 1219 1359 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03273 1092 1464 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03272 1359 2125 1092 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03271 2127 1464 1219 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03270 1217 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03269 2127 1215 1460 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03268 1215 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03267 2127 1222 1085 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03266 1085 1214 1215 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03265 1213 1211 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03264 2127 1981 1213 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03263 1064 1202 1199 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03262 2127 1196 1065 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03261 1061 1457 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03260 1199 1339 1061 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03259 1065 1198 1064 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03258 1063 1197 1065 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03257 1199 1849 1063 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03256 1194 1199 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03255 1202 1849 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03254 2127 1457 1196 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03253 1077 1884 1208 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03252 2127 1211 1077 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03251 1842 1208 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03250 1205 1842 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03249 1209 1610 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03248 2127 1211 1209 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03247 2127 1207 1453 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03246 1207 1753 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03245 2127 1204 1076 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03244 1076 1205 1207 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03243 1187 1190 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03242 1182 2126 1183 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03241 2127 1419 1182 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03240 2127 1191 1190 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03239 1192 1439 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03238 1192 1189 1191 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03237 1191 2125 1192 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03236 1428 2108 1188 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03235 1185 1183 1428 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03234 2127 1190 1188 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03233 1188 2105 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03232 1188 1184 1185 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03231 2127 1178 1179 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03230 1180 1291 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03229 1180 1177 1178 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03228 1178 2108 1180 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03227 1164 2101 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03226 2127 1174 1170 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03225 1173 1284 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03224 1173 1179 1174 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03223 1174 1175 1173 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03222 1172 2115 1175 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03221 2127 2058 1172 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03220 2127 1276 1162 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03219 1161 2105 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03218 1162 1187 1161 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03217 1424 1165 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03216 1169 1164 1166 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03215 1169 2108 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03214 2127 1168 1169 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03213 1166 1183 1165 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03212 1165 2105 1169 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03211 1236 1154 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03210 1158 1152 1155 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03209 1158 1884 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03208 2127 1891 1158 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03207 1155 1153 1154 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03206 1154 2058 1158 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03205 1146 1142 1145 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03204 2127 2108 1146 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03203 2127 1150 1151 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03202 1152 1151 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03201 2127 2115 1151 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03200 1151 1168 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03199 2127 1140 1153 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03198 1140 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03197 2127 1143 1144 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03196 1144 1145 1140 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03195 1143 1139 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03194 2127 1138 1139 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03193 1139 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03192 1119 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03191 2127 2108 1119 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03190 1280 1160 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03189 2127 1581 1160 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03188 1160 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03187 2127 1121 1629 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03186 1122 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03185 1122 1118 1121 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03184 1121 1119 1122 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03183 1113 1119 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03182 2127 1884 1113 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03181 1131 1126 1130 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03180 2127 1127 1133 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03179 1129 1541 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03178 1130 1128 1129 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03177 1133 1252 1131 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03176 1134 1261 1133 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03175 1130 1457 1134 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03174 1120 1130 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03173 1126 1457 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03172 2127 1541 1127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03171 1221 1097 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03170 2127 1099 1097 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03169 1097 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03168 2127 1096 1107 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03167 1107 1100 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03166 2127 1099 1100 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03165 1094 1096 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03164 1099 1101 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03163 2127 2113 1101 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03162 1101 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03161 1090 1086 1089 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03160 2127 1087 1093 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03159 1091 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03158 1089 1082 1091 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03157 1093 1226 1090 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03156 1088 1094 1093 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03155 1089 1884 1088 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03154 1620 1089 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03153 1086 1884 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03152 2127 2055 1087 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03151 1111 1105 1110 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03150 2127 1106 1109 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03149 1102 1753 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03148 1110 1170 1102 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03147 1109 1107 1111 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03146 1108 1346 1109 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03145 1110 2058 1108 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03144 1233 1110 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03143 1105 2058 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03142 2127 1753 1106 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03141 1073 1066 1072 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03140 2127 1067 1075 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03139 1070 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03138 1072 1068 1070 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03137 1075 1069 1073 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03136 1071 1213 1075 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03135 1072 1884 1071 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03134 1197 1072 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03133 1066 1884 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03132 2127 2055 1067 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03131 1211 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03130 2127 1081 1211 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03129 1084 2115 1083 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03128 2127 1081 1084 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03127 1470 1083 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03126 1060 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03125 2127 2122 1062 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03124 1069 1060 1059 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03123 1059 2122 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03122 1059 1062 1069 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03121 2127 2113 1059 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03120 2127 1074 1080 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03119 1080 1079 1081 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03118 1080 1078 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03117 1081 2122 1080 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03116 2127 1078 1079 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03115 1074 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03114 1184 1019 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03113 2127 1018 1019 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03112 1019 2126 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03111 2127 1006 1290 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03110 1290 1007 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03109 2127 2108 1007 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03108 916 1827 1177 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03107 2127 1419 916 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03106 929 1017 1015 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03105 2127 1012 930 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03104 924 1884 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03103 1015 1010 924 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03102 930 1009 929 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03101 931 1440 930 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03100 1015 2113 931 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03099 1254 1015 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03098 1017 2113 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03097 2127 1884 1012 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03096 898 989 990 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03095 2127 2108 898 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03094 1118 990 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03093 1003 1293 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03092 2127 1003 913 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03091 913 1004 1005 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03090 997 2088 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03089 2127 1000 1168 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03088 910 1004 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03087 910 1189 1000 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03086 1000 2126 910 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03085 1004 1001 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03084 2127 1018 1001 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03083 1001 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03082 908 1005 998 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03081 2127 2108 908 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03080 1276 998 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03079 903 1168 995 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03078 2127 2108 903 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03077 996 995 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03076 2127 997 1138 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03075 1138 991 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03074 2127 1273 991 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03073 987 986 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03072 2127 1006 986 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03071 986 984 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03070 904 1189 1273 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03069 2127 2125 904 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03068 1150 993 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03067 2127 2105 1150 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03066 1492 964 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03065 887 987 886 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03064 887 2123 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03063 2127 961 887 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_03062 886 970 964 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03061 964 962 887 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03060 962 960 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03059 2127 2058 960 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03058 960 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03057 2127 1273 969 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03056 970 969 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03055 2127 2108 969 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03054 969 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03053 2127 1113 974 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03052 974 971 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03051 974 2088 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03050 890 983 980 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03049 2127 977 895 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03048 891 1457 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03047 980 975 891 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03046 895 1651 890 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03045 894 979 895 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03044 980 1849 894 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03043 1128 980 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03042 983 1849 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03041 2127 1457 977 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_03040 971 948 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03039 2127 947 948 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03038 948 1956 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03037 961 1609 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03036 2105 2108 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03035 2127 956 1096 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03034 1096 958 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03033 2127 2113 958 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03032 950 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03031 2127 951 953 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03030 956 950 883 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03029 883 951 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03028 883 953 956 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03027 2127 2123 883 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03026 944 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03025 2127 2125 946 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03024 1078 944 877 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03023 877 2125 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03022 877 946 1078 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03021 2127 2108 877 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03020 1735 935 869 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03019 869 1753 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03018 868 2055 1735 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03017 2127 939 868 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03016 939 940 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_03015 2127 932 876 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03014 876 937 935 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03013 876 940 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03012 935 2108 876 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03011 2127 940 937 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03010 932 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03009 940 942 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03008 2127 2058 942 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03007 942 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03006 2127 1673 918 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03005 912 2123 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03004 918 911 912 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_03003 923 919 921 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03002 2127 917 922 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03001 915 2115 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_03000 921 914 915 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02999 922 918 923 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02998 920 1006 922 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02997 921 2105 920 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02996 1010 921 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02995 919 2105 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02994 2127 2115 917 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02993 2127 927 928 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02992 928 925 989 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02991 928 926 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02990 989 2123 928 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02989 2127 926 925 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02988 927 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02987 2127 909 914 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02986 863 989 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02985 864 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02984 865 2108 909 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02983 909 864 863 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02982 2127 1177 865 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02981 926 2126 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02980 2127 1898 926 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02979 907 1419 1006 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02978 2127 906 907 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02977 2127 902 1406 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02976 855 901 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02975 855 858 902 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02974 902 2105 855 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02973 862 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02972 2127 1005 862 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02971 1142 905 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02970 2127 2101 905 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02969 905 859 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02968 858 1419 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02967 2127 856 858 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02966 2127 1899 900 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02965 899 911 901 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02964 900 2105 899 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02963 2127 996 854 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02962 854 897 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02961 854 2093 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02960 853 984 896 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02959 2127 2113 853 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02958 897 896 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02957 889 888 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02956 2127 1827 888 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02955 888 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02954 984 889 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02953 852 889 892 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02952 852 1204 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02951 2127 1164 852 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02950 892 2058 852 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02949 893 892 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02948 884 1898 885 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02947 2127 2058 884 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02946 2127 849 979 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02945 979 850 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02944 2127 847 979 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02943 979 848 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02942 2127 2058 879 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02941 878 880 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02940 879 1280 878 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02939 881 1898 880 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02938 2127 1581 881 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02937 2127 885 850 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02936 850 846 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02935 850 984 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02934 845 2108 882 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02933 2127 2123 845 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02932 947 882 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02931 2127 2113 846 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02930 846 947 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02929 846 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02928 951 911 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02927 2127 2105 951 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02926 1654 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02925 2127 2108 1654 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02924 1609 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02923 2127 1753 1609 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02922 873 939 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02921 2127 873 875 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02920 875 951 874 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02919 2127 870 1082 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02918 872 871 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02917 1082 1884 872 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02916 1544 1541 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02915 2127 2113 840 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02914 840 2058 839 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02913 839 843 867 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02912 870 867 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02911 843 1078 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02910 742 2105 831 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02909 2127 835 742 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02908 830 831 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02907 743 834 836 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02906 743 2105 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02905 2127 835 743 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02904 836 2108 743 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02903 1009 836 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02902 740 1898 819 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02901 2127 1827 740 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02900 820 819 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02899 835 856 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02898 2127 1898 835 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02897 2127 826 1431 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02896 741 2115 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02895 741 830 826 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02894 826 824 741 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02893 818 820 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02892 2127 2105 818 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02891 805 820 736 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02890 736 2105 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02889 735 2108 805 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02888 2127 997 735 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02887 2127 809 1263 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02886 737 805 809 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02885 738 806 737 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02884 739 807 738 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02883 739 1162 2127 2127 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02882 2127 1884 739 2127 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02881 739 814 2127 2127 tp L=1U W=11U AS=22P AD=22P PS=26U PD=26U 
Mtr_02880 809 2058 739 2127 tp L=1U W=12U AS=24P AD=24P PS=28U PD=28U 
Mtr_02879 2127 862 814 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02878 814 818 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02877 814 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02876 734 820 803 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02875 2127 2108 734 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02874 802 803 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02873 2127 802 799 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02872 733 1142 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02871 799 2105 733 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02870 1827 773 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02869 2127 795 848 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02868 732 794 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02867 732 1884 795 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02866 795 859 732 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02865 2127 782 788 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02864 728 2113 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02863 788 802 728 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02862 785 792 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02861 730 854 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02860 2127 2058 730 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02859 730 1884 729 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02858 792 1753 731 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02857 729 788 730 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02856 729 2055 731 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02855 731 787 729 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02854 731 893 792 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02853 2127 773 769 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02852 770 769 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02851 2127 2105 769 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02850 769 766 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02849 2127 1138 782 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02848 727 856 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02847 782 780 727 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02846 2127 771 847 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02845 725 1884 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02844 847 770 725 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02843 773 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02842 2127 2123 773 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02841 726 1884 776 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02840 2127 782 726 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02839 849 776 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02838 1581 780 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02837 723 2055 759 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02836 2127 2122 723 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02835 780 745 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02834 2127 2113 745 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02833 745 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02832 761 1553 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02831 2127 759 761 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02830 751 747 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02829 2127 780 747 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02828 747 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02827 754 756 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02826 724 766 758 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02825 2127 2058 724 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02824 756 758 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02823 2127 2055 722 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02822 1214 755 722 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02821 722 756 1214 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02820 1346 750 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02819 2127 871 1346 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02818 2127 2055 752 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02817 721 754 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02816 752 751 721 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02815 911 926 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02814 834 720 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02813 2127 926 834 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02812 719 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02811 2127 1898 719 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02810 714 2105 715 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02809 2127 1293 714 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02808 716 715 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02807 717 718 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02806 718 1884 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02805 2127 2113 718 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02804 718 719 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02803 2127 1827 718 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02802 2127 709 1799 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02801 1799 708 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02800 1799 710 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02799 705 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02798 2127 715 705 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02797 707 715 706 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02796 2127 1142 707 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02795 708 706 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02794 2127 2108 712 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02793 712 2113 711 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02792 711 720 713 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02791 710 713 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02790 2127 2113 709 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02789 709 2088 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02788 709 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02787 704 843 703 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02786 2127 2122 704 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02785 701 703 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02784 2127 698 700 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02783 807 700 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02782 2127 2115 700 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02781 700 843 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02780 2127 697 794 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02779 794 699 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02778 2127 993 699 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02777 697 696 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02776 2127 2108 696 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02775 696 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02774 2127 799 702 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02773 702 705 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02772 702 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02771 694 785 695 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02770 694 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02769 2127 693 694 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02768 695 1849 694 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02767 692 695 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02766 2127 771 690 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02765 687 686 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02764 690 689 687 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02763 685 1898 771 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02762 2127 2055 685 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02761 2127 2113 688 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02760 689 856 688 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02759 688 2108 689 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02758 2127 691 693 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02757 693 690 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02756 2127 702 693 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02755 693 974 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02754 679 1899 678 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02753 2127 681 679 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02752 684 678 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02751 2127 1884 691 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02750 691 684 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02749 691 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02748 2127 676 677 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02747 675 1753 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02746 675 879 676 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02745 676 674 675 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02744 686 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02743 2127 683 686 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02742 680 2115 682 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02741 2127 1654 680 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02740 681 682 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02739 673 681 672 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02738 2127 2058 673 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02737 674 672 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02736 750 667 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02735 671 750 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02734 669 681 670 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02733 2127 1884 669 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02732 670 2058 671 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02731 668 670 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02730 667 666 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02729 2127 2113 666 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02728 666 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02727 755 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02726 2127 667 755 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02725 2127 664 871 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02724 871 665 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02723 2127 2113 665 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02722 856 650 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02721 552 2126 650 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02720 2127 2123 552 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02719 2127 1753 651 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02718 553 656 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02717 651 717 553 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02716 2127 659 554 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02715 656 1532 554 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02714 554 716 656 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02713 555 716 661 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02712 2127 2113 555 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02711 663 661 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02710 659 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02709 2127 2058 659 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02708 551 1164 636 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02707 2127 2108 551 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02706 638 636 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02705 649 2126 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02704 2127 1899 649 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02703 906 649 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02702 642 1673 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02701 2127 649 642 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02700 2127 642 641 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02699 806 641 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02698 2127 2113 641 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02697 641 638 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02696 2127 629 628 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02695 549 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02694 549 2115 629 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02693 629 1654 549 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02692 2127 701 550 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02691 634 2115 550 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02690 550 997 634 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02689 623 618 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02688 993 626 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02687 2127 997 626 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02686 626 623 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02685 2127 621 787 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02684 548 620 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02683 787 623 548 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02682 547 1899 618 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02681 2127 1164 547 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02680 2127 2105 621 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02679 621 612 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02678 2127 618 621 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02677 621 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02676 598 1654 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02675 2127 1898 598 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02674 2127 595 596 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02673 545 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02672 545 598 595 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02671 595 2058 545 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02670 546 600 603 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02669 546 598 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02668 2127 602 546 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02667 603 1849 546 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02666 975 603 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02665 602 611 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02664 611 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02663 2127 2123 611 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02662 611 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02661 2127 1764 611 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02660 543 2126 590 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02659 2127 588 543 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02658 2127 582 578 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02657 539 761 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02656 539 612 582 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02655 582 2058 539 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02654 2127 585 580 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02653 585 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02652 2127 1609 542 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02651 542 583 585 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02650 544 2113 592 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02649 2127 2125 544 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02648 612 592 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02647 2127 2122 541 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02646 540 590 589 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02645 541 1849 540 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02644 531 874 565 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02643 532 1544 531 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02642 533 1899 532 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02641 2127 560 533 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02640 2127 565 563 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02639 2127 563 534 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02638 566 752 534 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02637 534 589 566 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02636 2127 2122 579 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02635 538 2058 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02634 579 576 538 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02633 2127 572 567 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02632 572 566 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02631 2127 574 536 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02630 536 1457 572 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02629 557 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02628 2127 576 561 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02627 664 557 530 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02626 530 576 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02625 530 561 664 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02624 2127 2122 530 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02623 574 579 537 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02622 535 1753 574 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02621 2127 677 537 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02620 537 580 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02619 537 668 535 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02618 2127 527 528 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02617 529 528 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02616 2127 2113 528 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02615 528 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02614 517 663 516 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02613 2127 2058 517 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02612 2127 2058 523 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02611 524 522 523 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02610 523 663 524 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02609 520 2115 521 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02608 2127 519 520 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02607 522 521 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02606 518 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02605 2127 650 518 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02604 2127 1753 525 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02603 526 529 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02602 525 524 526 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02601 514 527 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02600 2127 514 513 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02599 513 1282 515 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02598 2127 2058 506 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02597 508 859 507 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02596 506 2108 508 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02595 511 2055 510 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02594 509 516 511 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02593 2127 1517 510 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02592 510 1884 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02591 510 515 509 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02590 2127 525 503 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02589 503 501 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02588 503 502 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02587 2127 1676 512 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02586 512 651 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02585 512 511 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02584 496 495 498 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02583 2127 1656 496 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02582 2127 499 497 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02581 500 494 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02580 500 628 499 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02579 499 1884 500 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02578 2127 493 501 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02577 493 491 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02576 2127 498 492 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02575 492 1884 493 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02574 490 503 489 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02573 490 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02572 2127 512 490 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02571 489 1849 490 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02570 488 489 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02569 504 1018 505 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02568 2127 2126 504 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02567 859 505 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02566 2127 476 600 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02565 600 477 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02564 600 497 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02563 2127 766 472 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02562 472 588 473 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02561 473 1753 471 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02560 491 471 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02559 2127 474 476 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02558 478 1884 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02557 476 634 478 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02556 486 483 485 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02555 2127 482 487 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02554 481 1541 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02553 485 479 481 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02552 487 488 486 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02551 484 692 487 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02550 485 1457 484 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02549 480 485 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02548 483 1457 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02547 2127 1541 482 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02546 475 1899 474 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02545 2127 2055 475 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02544 2127 461 463 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02543 462 469 464 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02542 463 465 462 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02541 465 466 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02540 2127 2105 466 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02539 466 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02538 470 2058 588 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02537 2127 2108 470 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02536 468 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02535 2127 2055 468 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02534 2127 612 469 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02533 469 467 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02532 2127 468 467 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02531 457 456 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02530 2127 2113 456 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02529 456 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02528 766 457 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02527 451 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02526 2127 453 455 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02525 452 451 454 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02524 454 453 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02523 454 455 452 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02522 2127 2122 454 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02521 460 465 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02520 2127 460 459 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02519 459 2058 1204 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02518 458 457 461 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02517 2127 2058 458 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02516 448 446 447 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02515 2127 444 449 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02514 445 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02513 447 443 445 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02512 449 452 448 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02511 450 1209 449 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02510 447 2058 450 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02509 1198 447 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02508 446 2058 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02507 2127 2055 444 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02506 502 1884 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02505 2127 434 502 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02504 2127 437 438 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02503 437 368 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02502 2127 519 367 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02501 367 2113 437 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02500 2127 433 434 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02499 434 438 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02498 434 518 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02497 368 527 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02496 370 1293 527 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02495 2127 2108 370 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02494 2127 429 433 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02493 433 2088 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02492 433 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02491 429 2123 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02490 2127 2105 429 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02489 2127 423 1419 2127 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_02488 1419 423 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02487 2127 1753 354 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02486 354 355 353 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02485 353 416 419 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02484 494 419 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02483 519 1164 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02482 2127 363 519 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02481 358 620 359 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02480 2127 1673 358 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02479 2127 2126 357 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02478 356 362 495 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02477 357 2115 356 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02476 2127 2105 361 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02475 361 2058 360 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02474 360 2115 424 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02473 620 424 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02472 362 429 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02471 416 415 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02470 2127 1464 415 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02469 415 2126 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02468 343 386 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02467 2127 474 343 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02466 2127 402 479 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02465 349 399 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02464 349 348 402 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02463 402 1457 349 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02462 2127 1899 342 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02461 341 1457 340 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02460 340 1764 345 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02459 342 396 341 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02458 396 394 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02457 2127 911 394 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02456 394 1581 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02455 2127 596 397 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02454 399 397 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02453 2127 390 397 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02452 397 345 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02451 407 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02450 2127 411 408 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02449 410 407 351 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02448 351 411 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02447 351 408 410 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02446 2127 2125 351 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02445 338 1884 387 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02444 2127 389 338 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02443 386 387 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02442 2127 1884 390 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02441 339 389 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02440 390 1898 339 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02439 352 1884 411 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02438 2127 1464 352 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02437 381 334 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02436 389 576 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02435 275 382 378 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02434 2127 376 276 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02433 271 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02432 378 377 271 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02431 276 410 275 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02430 274 381 276 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02429 378 2055 274 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02428 1538 378 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02427 382 2055 2127 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02426 2127 1764 376 2127 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_02425 333 2108 371 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02424 2127 2125 333 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02423 576 371 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02422 1757 1457 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02421 453 389 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02420 2127 2115 453 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02419 2127 332 330 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02418 331 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02417 331 1293 332 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02416 332 2108 331 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02415 2127 323 324 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02414 324 330 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02413 324 325 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02412 355 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02411 2127 1293 355 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02410 327 906 326 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02409 2127 2108 327 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02408 325 326 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02407 329 355 328 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02406 2127 2108 329 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02405 824 328 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02404 321 1753 322 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02403 2127 720 321 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02402 319 322 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02401 2127 1753 316 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02400 314 507 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02399 316 313 314 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02398 318 906 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02397 2127 1581 318 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02396 312 411 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02395 2127 312 311 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02394 311 310 313 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02393 2127 318 320 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02392 320 1884 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02391 320 1177 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02390 2127 320 317 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02389 317 315 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02388 2127 316 317 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02387 317 324 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02386 309 1899 308 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02385 2127 2122 309 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02384 305 306 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02383 2127 698 306 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02382 306 304 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02381 2127 302 301 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02380 303 319 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02379 303 1581 302 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02378 302 1884 303 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02377 1018 308 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02376 698 307 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02375 2127 308 307 2127 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_02374 304 294 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02373 2127 1884 294 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02372 294 583 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02371 292 1898 293 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02370 2127 304 292 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02369 291 293 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02368 2127 295 298 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02367 298 297 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02366 2127 301 298 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02365 298 343 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02364 2127 296 297 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02363 297 423 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02362 297 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02361 300 317 299 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02360 300 1764 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02359 2127 298 300 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02358 299 1849 300 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02357 348 299 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02356 2127 578 284 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02355 279 284 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02354 2127 280 284 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02353 284 290 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02352 287 289 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02351 2127 1753 289 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02350 289 386 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02349 2127 1764 290 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02348 288 291 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02347 290 287 288 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02346 2127 281 285 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02345 283 1899 282 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02344 282 1457 286 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02343 285 464 283 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02342 1764 1849 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02341 277 2115 278 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02340 2127 2058 277 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02339 272 278 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02338 273 272 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02337 2127 1753 270 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02336 560 270 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02335 2127 266 270 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02334 270 272 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02333 334 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02332 2127 2058 334 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02331 2127 1541 269 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02330 268 1899 267 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02329 267 1757 280 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02328 269 266 268 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02327 266 265 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02326 2127 911 265 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02325 265 334 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02324 1434 310 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02323 2127 720 1434 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02322 1673 230 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02321 233 1189 234 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02320 2127 2126 233 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02319 720 234 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02318 230 229 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02317 2127 2122 229 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02316 229 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02315 231 1898 232 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02314 2127 2123 231 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02313 1189 232 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02312 213 2105 215 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02311 2127 355 213 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02310 214 215 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02309 2127 2058 315 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02308 216 217 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02307 315 220 216 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02306 208 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02305 2127 2123 212 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02304 423 208 209 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02303 209 2123 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02302 209 212 423 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02301 2127 2122 209 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02300 217 214 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02299 221 226 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02298 226 230 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02297 2127 2105 226 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02296 226 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02295 2127 2058 226 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02294 2127 2108 219 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02293 220 310 219 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02292 219 1673 220 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02291 203 205 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02290 2127 203 204 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02289 204 1189 206 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02288 205 1581 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02287 2127 2126 205 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02286 2127 201 199 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02285 201 200 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02284 2127 1018 135 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02283 135 205 201 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02282 200 206 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02281 197 1673 198 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02280 2127 195 197 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02279 281 177 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02278 2127 198 177 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02277 177 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02276 125 1884 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02275 124 390 191 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02274 2127 1899 124 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02273 191 199 125 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02272 477 191 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02271 296 583 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02270 2127 1899 296 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02269 194 2126 196 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02268 2127 195 194 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02267 583 196 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02266 2127 2058 188 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02265 188 198 189 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02264 189 1899 190 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02263 295 190 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02262 179 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02261 2127 2126 179 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02260 2127 1884 183 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02259 184 186 183 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02258 183 683 184 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02257 186 1581 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02256 2127 1898 186 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02255 2127 174 235 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02254 111 279 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02253 111 182 174 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02252 174 1541 111 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02251 2127 2113 683 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02250 683 180 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02249 2127 179 180 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02248 2127 164 1068 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02247 106 162 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02246 106 168 164 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02245 164 2058 106 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02244 377 171 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02243 170 273 165 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02242 170 2055 2127 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02241 2127 169 170 2127 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_02240 165 167 171 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02239 171 1753 170 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02238 160 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02237 2127 2125 161 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02236 168 160 157 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02235 157 2125 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02234 157 161 168 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02233 2127 2113 157 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02232 173 168 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02231 162 272 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02230 152 2122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02229 2127 2055 152 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02228 1898 2122 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02227 2127 2122 1898 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02226 2127 2122 1898 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02225 1898 2122 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02224 2127 2113 148 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02223 148 1189 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02222 148 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02221 156 2105 155 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02220 2127 720 156 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02219 151 152 323 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02218 2127 195 151 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02217 1293 150 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02216 363 2108 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02215 2127 1899 363 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02214 2127 720 154 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02213 153 2108 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02212 154 310 153 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02211 149 363 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02210 2127 2125 147 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02209 147 2055 145 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02208 145 149 146 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02207 144 146 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02206 2127 2055 143 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02205 142 359 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02204 143 221 142 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02203 141 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02202 2127 362 141 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02201 2127 133 134 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02200 133 137 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02199 2127 1884 136 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02198 136 214 133 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02197 137 206 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02196 2127 140 138 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02195 139 144 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02194 139 141 140 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02193 140 2058 139 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02192 2127 150 128 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02191 128 127 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02190 2127 126 127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02189 2127 143 131 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02188 131 130 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02187 131 134 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02186 2127 128 130 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02185 130 138 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02184 130 129 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02183 123 122 129 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02182 2127 1764 123 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02181 132 1899 150 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02180 2127 2125 132 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02179 2127 453 122 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02178 122 121 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02177 2127 1898 121 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02176 116 390 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02175 2127 2055 117 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02174 118 184 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02173 117 119 118 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02172 2127 114 113 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02171 114 116 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02170 2127 179 115 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02169 115 2113 114 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02168 119 120 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02167 2127 1884 120 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02166 120 122 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02165 2127 107 169 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02164 108 2058 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02163 169 173 108 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02162 167 109 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02161 2127 110 109 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02160 109 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02159 443 107 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02158 2127 126 443 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02157 2127 110 126 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02156 126 112 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02155 2127 2058 112 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02154 103 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02153 2127 2108 104 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02152 110 103 105 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02151 105 2108 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02150 105 104 110 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02149 2127 2113 105 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02148 2127 310 69 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02147 69 68 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02146 2127 155 68 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02145 1753 2055 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02144 2127 2058 74 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02143 74 155 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02142 74 2113 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02141 10 1018 70 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02140 2127 2125 10 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02139 310 70 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02138 2127 77 71 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02137 71 74 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02136 71 310 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02135 2127 2108 12 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02134 12 2058 11 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02133 11 1018 78 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02132 77 78 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02131 2127 148 65 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02130 62 65 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02129 2127 69 65 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02128 65 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02127 2127 59 57 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02126 9 154 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02125 63 61 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02124 8 61 59 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02123 59 63 9 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02122 2127 69 8 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02121 7 2058 56 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02120 2127 2113 7 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02119 61 56 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02118 52 53 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02117 2127 1753 53 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02116 53 71 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02115 2127 50 49 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02114 50 2055 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02113 2127 305 5 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02112 5 62 50 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02111 6 1884 55 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02110 2127 2113 6 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02109 1282 55 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02108 195 42 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02107 2127 1764 48 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02106 4 49 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02105 48 52 4 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02104 2127 2055 44 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02103 44 1282 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02102 2127 42 44 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02101 44 1189 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02100 34 1457 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02099 2127 131 34 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02098 2127 272 41 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02097 41 40 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02096 2127 44 40 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02095 2127 36 182 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02094 182 31 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02093 2127 34 182 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02092 182 48 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02091 2127 57 36 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02090 36 41 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02089 36 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02088 23 22 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02087 2127 1898 22 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02086 22 2058 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02085 2127 117 27 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02084 27 24 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02083 27 1849 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02082 31 286 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02081 2127 27 31 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02080 2127 1753 24 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02079 3 23 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02078 24 113 3 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02077 1884 2058 2127 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02076 2127 18 107 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02075 107 14 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02074 2127 1884 14 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02073 2 2113 20 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02072 2127 2108 2 2127 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_02071 42 20 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02070 16 2125 2127 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02069 2127 42 17 2127 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02068 18 16 1 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02067 1 42 2127 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02066 1 17 18 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02065 2127 2125 1 2127 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_02064 2124 2123 2040 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02063 2044 2124 2120 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02062 2040 2122 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02061 2044 2125 2126 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02060 2126 2125 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02059 2044 2125 2126 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02058 2126 2125 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02057 2044 2120 2034 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02056 2034 2116 2119 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02055 2119 2117 2032 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02054 2032 2125 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02053 2044 2125 2116 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02052 2117 2120 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02051 2044 2120 2121 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02050 2044 2103 2101 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02049 2103 2102 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02048 2104 2107 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02047 2107 2111 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02046 2044 2105 2107 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02045 2044 2108 2018 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02044 2018 2111 2109 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02043 2044 2125 2025 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02042 2025 2110 2111 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02041 2111 2114 2024 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02040 2024 2123 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02039 2044 2123 2110 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02038 2114 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02037 2044 2093 1998 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02036 1998 2092 2095 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02035 2095 2113 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02034 2100 2102 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02033 2044 2123 2097 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02032 2005 2097 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02031 2098 2100 2005 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02030 2003 2123 2098 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02029 2044 2102 2003 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02028 2044 2095 2096 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02027 2044 2113 2115 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02026 2044 2122 2009 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02025 2009 2126 2102 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02024 2087 2122 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02023 2044 2126 2087 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02022 2044 2089 2088 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02021 2089 2087 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_02020 1979 2098 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02019 2044 2105 1979 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02018 1979 2108 2078 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02017 2078 2083 1979 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02016 2044 2078 2075 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02015 2080 2105 1983 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02014 1983 2083 2080 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02013 2044 2092 1983 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02012 2079 2080 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02011 2044 2087 1989 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02010 1989 2082 2083 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02009 2083 2084 1986 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02008 1986 2123 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02007 2044 2123 2082 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02006 2084 2087 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02005 2092 2090 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02004 2090 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02003 2044 2098 2090 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_02002 2044 2066 1965 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02001 1965 2065 2069 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_02000 2069 2067 1964 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01999 1964 2123 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01998 2044 2123 2065 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01997 2067 2066 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01996 2064 2113 1957 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01995 2044 2064 2063 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01994 1957 2069 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01993 2071 2113 1969 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01992 2044 2071 2070 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01991 1969 2075 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01990 2074 2072 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01989 2072 2075 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01988 2044 2115 2072 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01987 2054 2058 1943 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01986 2044 2054 2049 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01985 1943 2063 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01984 2044 2070 2046 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01983 2048 2046 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01982 2044 2058 2048 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01981 2044 2063 2052 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01980 2059 2052 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01979 2044 2058 2059 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01978 2057 2059 1952 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01977 1952 2062 2057 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01976 2044 2055 1952 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01975 2056 2057 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01974 2060 2058 1953 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01973 2044 2060 2062 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01972 1953 2070 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01971 2050 2048 1939 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01970 1939 2049 2050 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01969 2044 2055 1939 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01968 2045 2050 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01967 2043 2042 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01966 2042 2041 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01965 2044 2105 2042 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01964 2036 2035 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01963 2035 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01962 2044 2119 2035 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01961 2039 2037 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01960 2044 2115 2037 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01959 2038 2043 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01958 2037 2036 2038 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01957 2030 2033 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01956 2033 2119 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01955 2044 2105 2033 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01954 2028 2026 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01953 2044 2115 2026 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01952 2031 2030 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01951 2026 2029 2031 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01950 2017 2015 2016 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01949 2016 2113 2017 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01948 2044 2039 2016 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01947 2014 2017 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01946 2013 2109 2012 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01945 2044 2013 2011 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01944 2012 2010 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01943 2044 2019 2021 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01942 2021 2020 2022 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01941 2022 2027 2023 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01940 2023 2123 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01939 2044 2123 2020 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01938 2027 2019 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01937 2008 2104 2007 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01936 2044 2008 2015 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01935 2007 2010 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01934 2093 1997 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01933 1997 2022 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01932 2044 2105 1997 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01931 2044 1995 1987 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01930 1987 2092 1988 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01929 1988 2113 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01928 2044 2108 1996 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01927 1996 2022 1995 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01926 2044 2010 2004 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01925 2004 2000 2001 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01924 2001 2002 1999 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01923 1999 2122 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01922 2044 2122 2000 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01921 2002 2010 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01920 2010 2006 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01919 2006 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01918 2044 2126 2006 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01917 2044 2123 1993 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01916 1993 1990 1994 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01915 1994 1992 1991 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01914 1991 2108 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01913 2044 2108 1990 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01912 1992 2123 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01911 1974 1973 1975 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01910 1975 1976 1974 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01909 2044 2055 1975 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01908 1972 1974 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01907 1980 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01906 1982 2001 1981 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01905 2044 1980 1982 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01904 1977 1978 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01903 1978 2079 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01902 2044 2115 1978 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01901 2044 2074 1985 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01900 1984 1985 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01899 2044 1988 1984 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01898 1976 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01897 2044 2074 1976 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01896 1946 2058 1945 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01895 2044 1946 1947 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01894 1945 1966 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01893 1967 2122 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01892 2044 2108 1963 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01891 1961 1963 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01890 2066 1967 1961 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01889 1968 2108 2066 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01888 2044 2122 1968 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01887 1958 2055 1959 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01886 2044 1958 1956 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01885 1959 2113 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01884 1970 2113 1971 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01883 2044 1970 1966 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01882 1971 2079 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01881 2044 1966 1955 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01880 1954 1955 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01879 2044 2058 1954 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01878 2044 2066 1960 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01877 1962 1960 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01876 2044 2113 1962 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01875 2044 1935 1938 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01874 1940 1938 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01873 2044 2058 1940 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01872 2044 1934 1933 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01871 1934 1956 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01870 1950 1948 1951 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01869 1951 1954 1950 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01868 2044 2055 1951 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01867 1949 1950 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01866 1936 2058 1937 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01865 2044 1936 1948 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01864 1937 1935 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01863 1942 1940 1944 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01862 1944 1947 1942 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01861 2044 2055 1944 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01860 1941 1942 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01859 2044 1907 1837 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01858 1837 1908 2041 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01857 2041 1909 1836 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01856 1836 2125 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01855 2044 2125 1908 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01854 1909 1907 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01853 2044 1907 1900 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01852 2044 1902 1829 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01851 1829 2029 1903 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01850 1903 2115 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01849 2044 2108 1826 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01848 1826 1901 1902 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01847 2029 1906 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01846 1906 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01845 2044 2041 1906 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01844 1811 2113 1891 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01843 1891 2011 1811 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01842 1811 2028 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01841 1885 1887 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01840 2044 1884 1887 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01839 1804 1886 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01838 1887 2028 1804 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01837 1818 2113 1896 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01836 1896 1895 1818 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01835 1818 2039 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01834 2044 1899 1819 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01833 1819 1898 1907 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01832 1886 1889 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01831 2044 2113 1889 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01830 1806 2104 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01829 1889 1893 1806 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01828 1894 1893 1813 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01827 2044 1894 1895 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01826 1813 2109 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01825 2044 2123 1899 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01824 1899 2123 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01823 2044 2123 1899 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01822 1899 2123 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01821 2044 1885 1883 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01820 1877 1879 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01819 1879 1994 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01818 2044 2115 1879 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01817 2044 1878 1880 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01816 1798 2058 1881 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01815 1881 1880 1798 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01814 1798 1885 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01813 1973 1864 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01812 2044 1884 1973 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01811 2044 2096 1787 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01810 1787 1977 1878 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01809 2044 1988 1782 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01808 1782 2058 1871 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01807 2044 2058 1868 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01806 1871 1868 1781 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01805 1781 1872 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01804 1867 1871 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01803 2044 1873 1872 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01802 1873 1874 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01801 1874 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01800 2044 1994 1874 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01799 1866 2074 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01798 2044 1884 1866 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01797 1860 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01796 2044 1864 1860 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01795 1864 1857 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01794 1857 2069 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01793 2044 2115 1857 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01792 2044 2113 1756 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01791 1756 2058 1751 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01790 1751 1898 1855 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01789 1863 1866 1770 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01788 1770 1860 1863 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01787 2044 2055 1770 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01786 1858 1863 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01785 1850 1949 1748 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01784 1748 1853 1850 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01783 2044 1849 1748 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01782 1848 1850 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01781 2044 1855 1752 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01780 1752 1852 1853 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01779 1853 2055 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01778 2044 1852 1743 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01777 1743 1842 1843 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01776 1843 2055 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01775 1838 2113 1737 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01774 2044 1838 1935 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01773 1737 1899 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01772 1841 2045 1740 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01771 1740 1843 1841 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01770 2044 1849 1740 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01769 1839 1841 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01768 1847 2115 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01767 1847 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01766 2044 2058 1847 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01765 2044 1847 1852 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01764 2044 2115 1824 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01763 1824 1820 1823 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01762 1823 1821 1822 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01761 1825 1901 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01760 1731 2105 1821 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01759 2044 1825 1731 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01758 2044 2126 1828 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01757 1828 2121 1901 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01756 1901 1827 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01755 1831 1830 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01754 1830 2121 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01753 2044 2126 1830 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01752 1833 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01751 2044 2122 1832 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01750 1834 1832 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01749 2019 1833 1834 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01748 1835 2122 2019 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01747 2044 2125 1835 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01746 2044 1814 1816 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01745 1730 1822 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01744 1729 1817 1730 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01743 1814 1884 1729 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01742 1808 1807 1810 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01741 2044 1808 1812 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01740 1810 1809 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01739 1893 1803 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01738 1803 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01737 2044 1807 1803 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01736 1807 1805 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01735 1805 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01734 2044 1900 1805 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01733 1815 2108 1817 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01732 1817 1812 1815 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01731 1815 2104 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01730 2044 1797 1721 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01729 2044 1802 1725 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01728 1725 1883 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01727 1797 1753 1724 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01726 1724 1793 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01725 1725 2055 1797 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01724 1800 1799 1801 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01723 2044 1800 1802 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01722 1801 1884 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01721 1796 1794 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01720 2044 2113 1794 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01719 1720 2093 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01718 1794 1795 1720 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01717 1793 1790 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01716 2044 1791 1790 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01715 1718 1878 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01714 1790 2058 1718 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01713 1789 1788 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01712 2044 2113 1788 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01711 1716 1995 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01710 1788 1795 1716 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01709 2044 1884 1775 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01708 1773 2055 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01707 1777 1772 1778 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01706 1778 1884 1780 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01705 1780 1775 1779 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01704 1779 1776 1777 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01703 2044 2055 1777 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01702 1774 1773 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01701 1780 1784 1774 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01700 2044 1780 1762 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01699 2044 1796 1713 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01698 1713 2074 1714 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01697 1785 1981 1784 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01696 1784 1884 1785 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01695 1785 1783 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01694 1786 2126 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01693 1786 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01692 2044 2058 1786 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01691 2044 1786 1783 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01690 2044 1792 1791 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01689 2044 1796 1772 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01688 2044 1764 1765 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01687 1768 1763 1767 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01686 1767 1764 1769 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01685 1769 1765 1766 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01684 1766 1762 1768 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01683 2044 1757 1768 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01682 1760 1758 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01681 1769 1759 1760 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01680 1758 1757 2044 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01679 1761 1753 1763 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01678 1763 1754 1761 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01677 1761 1755 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01676 1746 1899 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01675 1746 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01674 2044 2058 1746 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01673 2044 1746 1749 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01672 1792 1771 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01671 1771 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01670 2044 1898 1771 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01669 1750 2096 1700 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01668 1700 1884 1750 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01667 2044 1749 1700 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01666 1754 1750 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01665 1741 1941 1694 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01664 1694 1745 1741 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01663 2044 1764 1694 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01662 1742 1741 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01661 2044 2122 1687 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01660 1687 2058 1747 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01659 2044 1744 1745 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01658 1693 1753 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01657 1697 2113 1693 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01656 1744 1747 1697 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01655 2044 1753 1736 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01654 1689 1736 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01653 2044 1747 1689 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01652 1738 1742 1691 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01651 1691 1839 1738 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01650 2044 1757 1691 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01649 1739 1738 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01648 1686 2108 1594 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01647 2044 1686 1685 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01646 1594 1684 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01645 2044 2036 1593 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01644 1593 1682 1683 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01643 1588 1674 1676 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01642 1676 1903 1588 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01641 1588 2058 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01640 2044 2108 1587 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01639 1587 1673 1820 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01638 2044 1679 1677 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01637 2044 1685 1591 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01636 1591 1678 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01635 1679 2115 1590 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01634 1590 1683 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01633 1591 2113 1679 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01632 2044 1795 1678 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01631 2044 2058 1666 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01630 1663 2055 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01629 1584 1677 1582 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01628 1582 2058 1667 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01627 1667 1666 1583 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01626 1583 1665 1584 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01625 2044 2055 1584 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01624 1580 1663 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01623 1667 1661 1580 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01622 2044 1667 1662 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01621 1795 1671 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01620 1671 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01619 2044 2111 1671 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01618 1578 2014 1661 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01617 1661 1884 1578 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01616 1578 1658 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01615 1658 1635 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01614 1635 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01613 2044 2126 1635 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01612 2044 1795 1568 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01611 1568 1654 1645 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01610 1645 2115 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01609 1576 2058 1657 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01608 1657 2014 1576 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01607 1576 1653 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01606 2044 1650 1651 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01605 2044 1816 1573 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01604 1573 1648 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01603 1650 1753 1574 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01602 1574 1881 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01601 1573 2055 1650 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01600 2044 1654 1575 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01599 1575 1893 1656 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01598 1656 2113 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01597 1647 1645 1571 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01596 1571 1656 1647 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01595 2044 2058 1571 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01594 1648 1647 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01593 2044 1632 1563 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01592 1563 1658 1634 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01591 1634 2055 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01590 1631 1972 1562 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01589 1562 1634 1631 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01588 2044 1849 1562 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01587 1628 1631 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01586 2044 1658 1638 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01585 2044 1629 1776 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01584 2044 1639 1637 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01583 2044 1642 1565 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01582 1565 1638 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01581 1639 2055 1564 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01580 1564 1657 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01579 1565 1753 1639 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01578 1643 2058 1566 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01577 2044 1643 1642 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01576 1566 1714 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01575 2044 1962 1552 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01574 1552 2058 1615 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01573 2044 2058 1617 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01572 1615 1617 1554 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01571 1554 1616 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01570 1624 1615 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01569 1612 1898 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01568 1612 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01567 2044 1609 1612 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01566 2044 1612 1755 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01565 1607 1977 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01564 2044 1884 1607 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01563 2044 2055 1625 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01562 1619 1764 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01561 1559 1867 1557 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01560 1557 2055 1621 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01559 1621 1625 1558 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01558 1558 1624 1559 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01557 2044 1764 1559 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01556 1556 1619 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01555 1621 1620 1556 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01554 2044 1621 1759 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01553 2044 1792 1608 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01552 2044 1962 1610 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01551 1598 1607 1543 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01550 1543 1596 1598 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01549 2044 2055 1543 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01548 1599 1598 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01547 1601 1599 1547 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01546 1547 1689 1601 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01545 2044 1764 1547 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01544 1603 1601 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01543 1605 1628 1549 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01542 1549 1603 1605 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01541 2044 1757 1549 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01540 1600 1605 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01539 1596 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01538 2044 1899 1596 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01537 2044 1684 1537 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01536 1532 1589 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01535 1589 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01534 2044 1831 1589 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01533 2044 1831 1534 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01532 1534 1533 1684 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01531 1674 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01530 2044 1577 1674 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01529 1592 1537 1536 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01528 1536 2108 1592 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01527 2044 1682 1536 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01526 1577 1592 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01525 2044 2109 1521 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01524 1524 1521 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01523 2044 1522 1524 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01522 1518 1577 1517 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01521 1517 2115 1518 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01520 1518 2096 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01519 1520 1581 1665 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01518 1665 2111 1520 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01517 1520 1579 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01516 1527 1585 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01515 2044 1529 1585 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01514 1526 1900 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01513 1585 2126 1526 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01512 1529 1586 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01511 1586 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01510 2044 2113 1586 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01509 2044 1581 1514 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01508 1514 1527 1515 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01507 1570 1572 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01506 2044 1884 1572 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01505 1503 1877 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01504 1572 1527 1503 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01503 1498 2058 1499 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01502 1499 1567 1498 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01501 1498 1570 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01500 2044 1884 1513 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01499 1507 2055 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01498 1512 1508 1509 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01497 1509 1884 1511 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01496 1511 1513 1510 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01495 1510 1515 1512 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01494 2044 2055 1512 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01493 1506 1507 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01492 1511 1504 1506 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01491 2044 1511 1505 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01490 1501 2058 1504 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01489 1504 1569 1501 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01488 1501 1570 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01487 2044 1473 1569 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01486 2044 1849 1494 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01485 1490 1757 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01484 1493 1721 1491 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01483 1491 1849 1496 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01482 1496 1494 1495 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01481 1495 1492 1493 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01480 2044 1757 1493 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01479 1489 1490 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01478 1496 1488 1489 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01477 2044 1496 1487 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01476 2044 1753 1484 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01475 1481 1849 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01474 1485 1479 1483 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01473 1483 1753 1482 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01472 1482 1484 1486 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01471 1486 1499 1485 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01470 2044 1849 1485 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01469 1480 1481 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01468 1482 1637 1480 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01467 2044 1482 1488 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01466 2044 1864 1472 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01465 1472 1629 1473 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01464 1560 1873 1478 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01463 2044 1560 1477 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01462 1478 1864 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01461 1479 1561 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01460 2044 1474 1561 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01459 1476 1473 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01458 1561 2058 1476 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01457 1632 1555 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01456 1555 1470 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01455 2044 1884 1555 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01454 2044 1464 1616 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01453 2044 1632 1468 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01452 1468 1553 1469 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01451 1469 2055 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01450 1551 1858 1466 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01449 1466 1469 1551 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01448 2044 1764 1466 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01447 1463 1551 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01446 1550 1463 1462 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01445 1462 1460 1550 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01444 2044 1457 1462 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01443 1546 1550 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01442 2044 1769 1448 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01441 1448 1539 1447 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01440 1447 1540 1446 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01439 1545 2056 1455 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01438 1455 1453 1545 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01437 2044 1764 1455 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01436 1456 1545 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01435 1450 1542 1540 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01434 1540 1739 1450 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01433 1450 1541 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01432 1548 1848 1459 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01431 1459 1456 1548 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01430 2044 1457 1459 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01429 1542 1548 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01428 1452 1546 1539 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01427 1539 1600 1452 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01426 1452 1544 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01425 2044 1441 1337 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01424 1337 2108 1444 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01423 2044 2108 1445 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01422 1444 1445 1336 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01421 1336 2019 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01420 1440 1444 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01419 2044 1439 1533 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01418 1433 1435 1332 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01417 1332 2113 1433 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01416 2044 1431 1332 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01415 1567 1433 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01414 1333 2108 1435 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01413 1435 1438 1334 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01412 2044 1434 1333 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01411 1334 1522 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01410 2044 2108 1438 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01409 2044 1533 1335 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01408 1335 1673 1441 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01407 2044 1428 1429 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01406 2044 2115 1422 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01405 1423 1884 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01404 1331 1424 1330 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01403 1330 2115 1427 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01402 1427 1422 1329 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01401 1329 1429 1331 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01400 2044 1884 1331 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01399 1328 1423 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01398 1427 1896 1328 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01397 2044 1427 1420 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01396 2044 2105 1412 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01395 1413 2113 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01394 1324 1417 1323 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01393 1323 2105 1415 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01392 1415 1412 1322 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01391 1322 1900 1324 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01390 2044 2113 1324 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01389 1321 1413 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01388 1415 1406 1321 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01387 2044 1415 1508 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01386 2044 1673 1325 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01385 1325 1899 1417 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01384 2044 1809 1327 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01383 1327 2101 1522 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01382 2044 2125 1326 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01381 1326 1419 1809 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01380 2044 2055 1382 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01379 1383 1849 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01378 1314 1420 1313 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01377 1313 2055 1386 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01376 1386 1382 1312 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01375 1312 1384 1314 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01374 2044 1849 1314 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01373 1311 1383 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01372 1386 1394 1311 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01371 2044 1386 1378 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01370 2044 1714 1407 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01369 2044 2058 1396 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01368 1397 2055 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01367 1319 1395 1318 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01366 1318 2058 1402 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01365 1402 1396 1320 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01364 1320 1401 1319 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01363 2044 2055 1319 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01362 1317 1397 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01361 1402 1398 1317 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01360 2044 1402 1394 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01359 2044 1877 1316 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01358 1316 1464 1401 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01357 1315 1567 1393 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01356 1393 1884 1315 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01355 1315 1391 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01354 1310 1884 1384 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01353 1384 1984 1310 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01352 1310 1373 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01351 2044 1391 1474 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01350 1553 1368 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01349 1368 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01348 2044 2105 1368 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01347 1309 1477 1398 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01346 1398 1884 1309 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01345 1309 1553 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01344 1366 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01343 1308 1365 1391 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01342 2044 1366 1308 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01341 1358 1361 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01340 2044 1360 1361 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01339 1305 1359 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01338 1361 2058 1305 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01337 1364 2058 1306 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01336 2044 1364 1363 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01335 1306 1365 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01334 2044 1470 1307 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01333 1307 1981 1365 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01332 2044 1553 1360 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01331 1464 1375 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01330 1375 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01329 2044 2105 1375 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01328 2044 1609 1355 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01327 1349 1347 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01326 2044 1351 1347 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01325 1301 1346 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01324 1347 2058 1301 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01323 1373 1356 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01322 2044 2058 1356 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01321 1304 1470 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01320 1356 1610 1304 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01319 2044 1753 1341 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01318 1338 1849 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01317 1299 1358 1300 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01316 1300 1753 1343 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01315 1343 1341 1298 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01314 1298 1349 1299 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01313 2044 1849 1299 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01312 1297 1338 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01311 1343 1350 1297 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01310 2044 1343 1339 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01309 2044 1352 1350 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01308 2044 1363 1303 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01307 1303 1608 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01306 1352 2125 1302 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01305 1302 1355 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01304 1303 2055 1352 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01303 2044 1373 1351 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01302 1289 2105 1288 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01301 1288 1434 1289 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01300 1289 1290 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01299 2044 1290 1291 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01298 1281 1884 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01297 2044 1428 1281 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01296 1682 1295 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01295 2044 2105 1295 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01294 1296 1294 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01293 1295 1293 1296 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01292 2044 2125 1292 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01291 1292 1900 1294 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01290 1439 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01289 2044 1419 1439 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01288 2044 1431 1287 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01287 1395 1285 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01286 2044 1287 1285 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01285 1286 1288 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01284 1285 2115 1286 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01283 1277 1275 1653 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01282 1653 1279 1277 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01281 1277 1281 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01280 2044 1282 1283 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01279 1283 1900 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01278 1284 1524 1283 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01277 1283 2113 1284 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01276 2044 1276 1278 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01275 1278 2115 1279 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01274 2044 1280 1579 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01273 1271 2058 1270 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01272 1270 1407 1271 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01271 1271 1653 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01270 2044 2055 1269 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01269 1264 1849 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01268 1266 1263 1268 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01267 1268 2055 1267 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01266 1267 1269 1265 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01265 1265 1270 1266 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01264 2044 1849 1266 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01263 1262 1264 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01262 1267 1662 1262 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01261 2044 1267 1261 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01260 1272 1273 1274 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01259 1274 1827 1272 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01258 2044 2108 1274 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01257 1275 1272 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01256 2044 2055 1260 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01255 1255 1764 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01254 1256 1254 1257 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01253 1257 2055 1259 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01252 1259 1260 1258 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01251 1258 1393 1256 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01250 2044 1764 1256 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01249 1253 1255 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01248 1259 1505 1253 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01247 2044 1259 1252 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01246 2044 1757 1249 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01245 1245 1541 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01244 1251 1378 1250 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01243 1250 1757 1247 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01242 1247 1249 1248 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01241 1248 1246 1251 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01240 2044 1541 1251 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01239 1244 1245 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01238 1247 1487 1244 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01237 2044 1247 1243 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01236 2044 1789 1227 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01235 1227 1977 1228 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01234 2044 1228 1232 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01233 1232 2058 1231 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01232 2044 2058 1229 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01231 1231 1229 1230 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01230 1230 1359 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01229 1235 1231 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01228 2044 1789 1226 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01227 2044 2055 1239 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01226 1237 1764 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01225 1240 1236 1242 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01224 1242 2055 1241 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01223 1241 1239 1238 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01222 1238 1235 1240 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01221 2044 1764 1240 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01220 1234 1237 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01219 1241 1233 1234 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01218 2044 1241 1246 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01217 1225 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01216 2044 1977 1225 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01215 1223 1221 1224 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01214 1224 1225 1223 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01213 2044 2055 1224 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01212 1222 1223 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01211 2044 1464 1220 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01210 1220 1217 1359 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01209 1359 1219 1218 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01208 1218 2125 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01207 2044 2125 1217 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01206 1219 1464 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01205 1215 1222 1216 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01204 1216 1214 1215 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01203 2044 1849 1216 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01202 1460 1215 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01201 2044 1211 1212 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01200 1212 1981 1213 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01199 2044 1849 1202 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01198 1196 1457 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01197 1201 1198 1203 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01196 1203 1849 1199 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01195 1199 1202 1200 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01194 1200 1197 1201 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01193 2044 1457 1201 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01192 1195 1196 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01191 1199 1339 1195 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01190 2044 1199 1194 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01189 1842 1208 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01188 1208 1211 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01187 2044 1884 1208 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01186 2044 1842 1205 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01185 2044 1610 1210 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01184 1210 1211 1209 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01183 1207 1204 1206 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01182 1206 1205 1207 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01181 2044 1753 1206 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01180 1453 1207 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01179 2044 1190 1187 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01178 1183 1419 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01177 2044 2126 1183 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01176 1190 1191 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01175 2044 1439 1191 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01174 1058 1189 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01173 1191 2125 1058 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01172 1056 1184 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01171 1057 1190 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01170 2044 1183 1056 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01169 1056 2108 1428 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01168 1428 2105 1057 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01167 1179 1178 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01166 2044 1291 1178 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01165 1055 1177 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01164 1178 2108 1055 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01163 2044 2101 1164 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01162 1170 1174 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01161 2044 1284 1174 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01160 1054 1179 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01159 1174 1175 1054 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01158 1175 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01157 2044 2115 1175 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01156 1051 2105 1162 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01155 1162 1187 1051 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01154 1051 1276 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01153 2044 1165 1424 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01152 2044 1183 1052 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01151 1052 1164 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01150 1165 2108 1053 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01149 1053 1168 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01148 1052 2105 1165 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01147 2044 1154 1236 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01146 2044 1153 1048 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01145 1048 1152 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01144 1154 1884 1049 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01143 1049 1891 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_01142 1048 2058 1154 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01141 1145 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01140 2044 1142 1145 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01139 2044 1151 1152 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01138 1046 1150 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01137 1047 1168 1046 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01136 1151 2115 1047 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01135 1140 1143 1045 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01134 1045 1145 1140 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01133 2044 2113 1045 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01132 1153 1140 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01131 1139 2108 1044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01130 2044 1139 1143 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01129 1044 1138 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01128 2044 2123 1039 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01127 1039 2108 1119 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01126 1160 2125 1050 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01125 2044 1160 1280 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01124 1050 1581 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01123 1629 1121 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01122 2044 2113 1121 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01121 1040 1118 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01120 1121 1119 1040 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01119 2044 1119 1038 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01118 1038 1884 1113 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01117 2044 1457 1126 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01116 1127 1541 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01115 1042 1252 1041 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01114 1041 1457 1130 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01113 1130 1126 1043 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01112 1043 1261 1042 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01111 2044 1541 1042 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01110 988 1127 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01109 1130 1128 988 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01108 2044 1130 1120 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01107 1097 2058 1032 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01106 2044 1097 1221 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01105 1032 1099 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01104 1100 1099 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01103 1033 1096 1107 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01102 2044 1100 1033 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01101 2044 1096 1094 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01100 1101 2123 1034 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01099 2044 1101 1099 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01098 1034 2113 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01097 2044 1884 1086 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01096 1087 2055 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01095 1031 1226 1029 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01094 1029 1884 1089 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01093 1089 1086 1030 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01092 1030 1094 1031 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01091 2044 2055 1031 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01090 955 1087 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01089 1089 1082 955 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01088 2044 1089 1620 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01087 2044 2058 1105 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01086 1106 1753 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01085 1036 1107 1035 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01084 1035 2058 1110 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01083 1110 1105 1037 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01082 1037 1346 1036 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01081 2044 1753 1036 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01080 966 1106 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01079 1110 1170 966 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01078 2044 1110 1233 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01077 2044 1884 1066 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01076 1067 2055 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01075 1025 1069 1024 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01074 1024 1884 1072 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01073 1072 1066 1023 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01072 1023 1213 1025 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01071 2044 2055 1025 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01070 938 1067 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01069 1072 1068 938 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01068 2044 1072 1197 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01067 2044 2113 1028 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01066 1028 1081 1211 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01065 1470 1083 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01064 1083 1081 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01063 2044 2115 1083 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01062 1062 2122 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01061 2044 2113 1060 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01060 1022 1060 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01059 1069 1062 1022 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01058 1021 2113 1069 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01057 2044 2122 1021 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01056 2044 1078 1026 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01055 1026 1074 1081 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01054 1081 1079 1027 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01053 1027 2122 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01052 2044 2122 1074 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01051 1079 1078 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01050 1019 2126 1020 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01049 2044 1019 1184 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01048 1020 1018 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01047 1007 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01046 1008 1006 1290 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01045 2044 1007 1008 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01044 1177 1419 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01043 2044 1827 1177 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01042 2044 2113 1017 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_01041 1012 1884 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_01040 1014 1009 1013 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01039 1013 2113 1015 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01038 1015 1017 1016 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01037 1016 1440 1014 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01036 2044 1884 1014 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01035 1011 1012 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01034 1015 1010 1011 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01033 2044 1015 1254 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01032 1118 990 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01031 990 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01030 2044 989 990 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01029 2044 1293 1003 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01028 1005 1003 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01027 2044 1004 1005 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01026 2044 2088 997 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01025 1168 1000 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01024 2044 1004 1000 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01023 999 1189 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01022 1000 2126 999 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01021 1001 2125 1002 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01020 2044 1001 1004 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01019 1002 1018 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01018 1276 998 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01017 998 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01016 2044 1005 998 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01015 996 995 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01014 995 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01013 2044 1168 995 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01012 991 1273 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01011 992 997 1138 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01010 2044 991 992 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01009 986 984 985 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01008 2044 986 987 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01007 985 1006 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01006 1273 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01005 2044 1189 1273 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_01004 2044 993 994 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01003 994 2105 1150 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01002 2044 964 1492 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01001 2044 970 965 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01000 965 987 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00999 964 2123 963 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00998 963 961 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00997 965 962 964 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00996 960 2055 959 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00995 2044 960 962 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00994 959 2058 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00993 2044 969 970 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00992 967 1273 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00991 968 2113 967 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00990 969 2108 968 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00989 2044 2088 973 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00988 973 1113 972 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00987 972 971 974 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00986 2044 1849 983 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00985 977 1457 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00984 982 1651 978 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00983 978 1849 980 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00982 980 983 981 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00981 981 979 982 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00980 2044 1457 982 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00979 976 977 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00978 980 975 976 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00977 2044 980 1128 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00976 948 1956 949 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00975 2044 948 971 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00974 949 947 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00973 2044 1609 961 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00972 2044 2108 2105 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00971 958 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00970 957 956 1096 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00969 2044 958 957 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00968 953 951 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00967 2044 2123 950 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00966 954 950 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00965 956 953 954 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00964 952 2123 956 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00963 2044 951 952 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00962 946 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00961 2044 2108 944 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00960 945 944 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00959 1078 946 945 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00958 943 2108 1078 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00957 2044 2125 943 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00956 2044 939 933 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00955 933 2055 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00954 1735 935 933 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00953 933 1753 1735 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00952 2044 940 939 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00951 2044 940 936 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00950 936 932 935 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00949 935 937 934 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00948 934 2108 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00947 2044 2108 932 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00946 937 940 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00945 942 2113 941 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00944 2044 942 940 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00943 941 2058 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00942 821 2123 918 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00941 918 911 821 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00940 821 1673 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00939 2044 2105 919 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00938 917 2115 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00937 827 918 828 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00936 828 2105 921 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00935 921 919 829 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00934 829 1006 827 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00933 2044 2115 827 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00932 823 917 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00931 921 914 823 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00930 2044 921 1010 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00929 2044 926 833 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00928 833 927 989 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00927 989 925 832 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00926 832 2123 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00925 2044 2123 927 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00924 925 926 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00923 2044 989 815 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00922 815 2108 909 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00921 2044 2108 864 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00920 909 864 816 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00919 816 1177 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00918 914 909 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00917 2044 2126 866 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00916 866 1898 926 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00915 1006 906 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00914 2044 1419 1006 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00913 1406 902 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00912 2044 901 902 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00911 801 858 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00910 902 2105 801 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00909 2044 2108 861 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00908 861 1005 862 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00907 905 859 860 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00906 2044 905 1142 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00905 860 2101 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00904 2044 1419 857 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00903 857 856 858 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00902 2044 2105 901 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00901 901 1899 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00900 901 911 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00899 2044 2093 797 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00898 797 996 798 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00897 798 897 854 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00896 897 896 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00895 896 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00894 2044 984 896 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00893 888 2108 851 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00892 2044 888 889 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00891 851 1827 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00890 2044 889 984 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00889 790 889 892 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00888 2044 2058 790 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00887 786 1204 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00886 892 1164 786 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00885 2044 892 893 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00884 885 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00883 2044 1898 885 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00882 2044 848 778 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00881 778 849 777 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00880 777 850 779 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00879 779 847 979 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00878 762 880 879 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00877 879 1280 762 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00876 762 2058 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00875 880 1581 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00874 2044 1898 880 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00873 2044 984 775 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00872 775 885 774 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00871 774 846 850 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00870 947 882 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00869 882 2123 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00868 2044 2108 882 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00867 2044 2125 767 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00866 767 2113 765 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00865 765 947 846 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00864 2044 911 842 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00863 842 2105 951 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00862 2044 2125 844 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00861 844 2108 1654 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00860 2044 2058 841 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00859 841 1753 1609 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00858 2044 939 873 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00857 874 873 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00856 2044 951 874 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00855 749 871 1082 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00854 1082 1884 749 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00853 749 870 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00852 2044 1541 1544 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00851 867 843 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00850 867 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00849 2044 2058 867 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00848 2044 867 870 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00847 2044 1078 843 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00846 830 831 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00845 831 835 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00844 2044 2105 831 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00843 837 834 836 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00842 2044 2108 837 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00841 838 2105 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00840 836 835 838 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00839 2044 836 1009 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00838 820 819 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00837 819 1827 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00836 2044 1898 819 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00835 2044 856 822 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00834 822 1898 835 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00833 1431 826 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00832 2044 2115 826 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00831 825 830 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00830 826 824 825 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00829 2044 820 817 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00828 817 2105 818 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00827 2044 997 804 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00826 804 2108 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00825 805 820 804 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00824 804 2105 805 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00823 1263 809 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00822 808 2058 809 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00821 2044 805 808 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00820 808 806 2044 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00819 2044 807 808 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00818 809 814 811 2044 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_00817 811 1884 810 2044 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_00816 810 1162 2044 2044 tn L=1U W=8U AS=16P AD=16P PS=20U PD=20U 
Mtr_00815 2044 2113 812 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00814 812 862 813 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00813 813 818 814 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00812 802 803 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00811 803 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00810 2044 820 803 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00809 800 1142 799 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00808 799 2105 800 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00807 800 802 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00806 2044 773 1827 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00805 848 795 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00804 2044 794 795 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00803 796 1884 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00802 795 859 796 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00801 783 2113 788 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00800 788 802 783 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00799 783 782 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00798 791 787 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00797 2044 788 789 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00796 784 854 792 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00795 2044 2058 784 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00794 785 792 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00793 792 2055 791 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00792 789 1884 792 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00791 792 893 793 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00790 793 1753 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00789 2044 769 770 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00788 764 773 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00787 768 766 764 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00786 769 2105 768 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00785 781 856 782 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00784 782 780 781 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00783 781 1138 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00782 772 1884 847 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00781 847 770 772 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00780 772 771 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00779 2044 2125 763 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00778 763 2123 773 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00777 849 776 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00776 776 782 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00775 2044 1884 776 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00774 2044 780 1581 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00773 759 2122 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00772 2044 2055 759 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00771 745 2108 744 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00770 2044 745 780 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00769 744 2113 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00768 2044 1553 760 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00767 760 759 761 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00766 747 2058 748 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00765 2044 747 751 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00764 748 780 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00763 2044 756 754 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00762 756 758 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00761 758 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00760 2044 766 758 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00759 2044 755 757 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00758 757 756 1214 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00757 1214 2055 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00756 2044 750 746 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00755 746 871 1346 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00754 753 754 752 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00753 752 751 753 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00752 753 2055 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00751 2044 926 911 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00750 2044 720 662 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00749 662 926 834 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00748 2044 2108 657 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00747 657 1898 719 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00746 715 1293 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00745 2044 2105 715 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00744 2044 715 716 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00743 654 719 653 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00742 2044 1884 658 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00741 653 1827 718 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00740 658 2113 654 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00739 2044 718 717 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00738 2044 710 645 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00737 645 709 643 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00736 643 708 1799 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00735 2044 2113 637 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00734 637 715 705 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00733 708 706 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00732 706 1142 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00731 2044 715 706 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00730 713 720 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00729 713 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00728 2044 2113 713 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00727 2044 713 710 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00726 2044 2108 647 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00725 647 2113 646 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00724 646 2088 709 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00723 701 703 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00722 703 2122 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00721 2044 843 703 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00720 2044 700 807 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00719 625 698 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00718 630 843 625 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00717 700 2115 630 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00716 699 993 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00715 622 697 794 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00714 2044 699 622 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00713 696 2055 619 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00712 2044 696 697 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00711 619 2108 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00710 2044 2058 633 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00709 633 799 631 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00708 631 705 702 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00707 617 785 695 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00706 2044 1849 617 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00705 616 1764 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00704 695 693 616 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00703 2044 695 692 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00702 597 686 690 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00701 690 689 597 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00700 597 771 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00699 771 2055 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00698 2044 1898 771 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00697 2044 856 599 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00696 599 2108 689 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00695 689 2113 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00694 2044 974 605 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00693 605 691 607 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00692 607 690 606 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00691 606 702 693 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00690 684 678 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00689 678 681 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00688 2044 1899 678 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00687 2044 2122 587 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00686 587 1884 586 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00685 586 684 691 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00684 677 676 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00683 2044 1753 676 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00682 575 879 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00681 676 674 575 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00680 2044 2058 591 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00679 591 683 686 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00678 681 682 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00677 682 1654 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00676 2044 2115 682 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00675 674 672 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00674 672 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00673 2044 681 672 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00672 2044 667 750 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00671 570 681 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00670 2044 1884 570 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00669 570 750 670 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00668 670 2058 570 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00667 2044 670 668 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00666 666 2122 562 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00665 2044 666 667 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00664 562 2113 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00663 2044 2058 564 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00662 564 667 755 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00661 665 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00660 559 664 871 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00659 2044 665 559 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00658 2044 650 856 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00657 650 2123 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00656 2044 2126 650 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00655 652 656 651 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00654 651 717 652 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00653 652 1753 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00652 2044 1532 655 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00651 655 716 656 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00650 656 659 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00649 663 661 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00648 661 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00647 2044 716 661 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00646 2044 2113 660 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00645 660 2058 659 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00644 638 636 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00643 636 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00642 2044 1164 636 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00641 2044 2126 648 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00640 648 1899 649 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00639 2044 649 906 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00638 2044 1673 644 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00637 644 649 642 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00636 2044 641 806 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00635 639 642 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00634 640 638 639 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00633 641 2113 640 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00632 628 629 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00631 2044 2123 629 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00630 632 2115 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00629 629 1654 632 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00628 2044 2115 635 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00627 635 997 634 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00626 634 701 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00625 2044 618 623 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00624 626 623 627 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00623 2044 626 993 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00622 627 997 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00621 624 620 787 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00620 787 623 624 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00619 624 621 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00618 618 1164 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00617 2044 1899 618 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00616 2044 2058 615 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00615 615 2105 613 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00614 613 612 614 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00613 614 618 621 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00612 2044 1654 593 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00611 593 1898 598 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00610 596 595 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00609 2044 2055 595 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00608 594 598 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00607 595 2058 594 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00606 604 600 603 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00605 2044 1849 604 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00604 601 598 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00603 603 602 601 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00602 2044 603 975 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00601 609 2058 608 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00600 2044 2055 610 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00599 608 1764 611 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00598 610 2123 609 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00597 2044 611 602 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00596 590 588 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00595 2044 2126 590 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00594 578 582 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00593 2044 761 582 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00592 581 612 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00591 582 2058 581 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00590 585 1609 584 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00589 584 583 585 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00588 2044 1764 584 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00587 580 585 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00586 612 592 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00585 592 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00584 2044 2113 592 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00583 2044 1849 589 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00582 589 2122 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00581 589 590 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00580 565 560 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00579 2044 874 565 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00578 2044 1899 565 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00577 565 1544 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00576 563 565 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00575 2044 752 568 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00574 568 589 566 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00573 566 563 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00572 577 2058 579 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00571 579 576 577 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00570 577 2122 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00569 572 574 571 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00568 571 1457 572 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00567 2044 566 571 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00566 567 572 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00565 561 576 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00564 2044 2122 557 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00563 558 557 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00562 664 561 558 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00561 556 2122 664 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00560 2044 576 556 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00559 569 668 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00558 573 677 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00557 2044 1753 569 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00556 569 579 574 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00555 574 580 573 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00554 2044 528 529 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00553 441 527 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00552 442 2058 441 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00551 528 2113 442 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00550 516 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00549 2044 663 516 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00548 2044 522 439 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00547 439 663 524 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00546 524 2058 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00545 522 521 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00544 521 519 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00543 2044 2115 521 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00542 2044 2108 432 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00541 432 650 518 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00540 440 529 525 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00539 525 524 440 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00538 440 1753 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00537 2044 527 514 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00536 515 514 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00535 2044 1282 515 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00534 2044 2108 507 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00533 507 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00532 507 859 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00531 426 515 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00530 425 1517 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00529 2044 516 426 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00528 426 2055 511 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00527 511 1884 425 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00526 2044 502 421 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00525 421 525 422 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00524 422 501 503 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00523 2044 511 428 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00522 428 1676 427 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00521 427 651 512 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00520 498 1656 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00519 2044 495 498 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00518 497 499 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00517 2044 494 499 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00516 420 628 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00515 499 1884 420 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00514 493 498 417 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00513 417 1884 493 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00512 2044 491 417 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00511 501 493 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00510 414 503 489 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00509 2044 1849 414 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00508 412 1764 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00507 489 512 412 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00506 2044 489 488 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00505 859 505 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00504 505 2126 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00503 2044 1018 505 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00502 2044 497 401 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00501 401 476 400 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00500 400 477 600 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00499 471 1753 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00498 471 766 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00497 2044 588 471 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00496 2044 471 491 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00495 398 1884 476 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00494 476 634 398 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00493 398 474 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00492 2044 1457 483 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00491 482 1541 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00490 405 488 406 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00489 406 1457 485 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00488 485 483 404 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00487 404 692 405 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00486 2044 1541 405 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00485 403 482 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00484 485 479 403 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00483 2044 485 480 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00482 474 2055 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00481 2044 1899 474 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00480 2044 465 464 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00479 464 461 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00478 464 469 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00477 466 2113 388 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00476 2044 466 465 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00475 388 2105 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00474 588 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00473 2044 2058 588 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00472 2044 2122 393 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00471 393 2055 468 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00470 467 468 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00469 392 612 469 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00468 2044 467 392 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00467 456 2125 385 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00466 2044 456 457 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00465 385 2113 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00464 2044 457 766 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00463 455 453 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00462 2044 2122 451 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00461 380 451 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00460 452 455 380 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00459 384 2122 452 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00458 2044 453 384 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00457 2044 465 460 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00456 1204 460 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00455 2044 2058 1204 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00454 461 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00453 2044 457 461 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00452 2044 2058 446 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00451 444 2055 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00450 373 452 374 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00449 374 2058 447 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00448 447 446 375 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00447 375 1209 373 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00446 2044 2055 373 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00445 372 444 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00444 447 443 372 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00443 2044 447 1198 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00442 2044 1884 366 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00441 366 434 502 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00440 437 519 369 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00439 369 2113 437 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00438 2044 368 369 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00437 438 437 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00436 2044 518 436 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00435 436 433 435 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00434 435 438 434 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00433 2044 527 368 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00432 527 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00431 2044 1293 527 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00430 2044 2113 430 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00429 430 429 431 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00428 431 2088 433 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00427 2044 2123 365 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00426 365 2105 429 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00425 2044 423 1419 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00424 1419 423 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00423 419 416 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00422 419 1753 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00421 2044 355 419 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00420 2044 419 494 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00419 2044 1164 364 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00418 364 363 519 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00417 359 1673 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00416 2044 620 359 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00415 2044 2115 495 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00414 495 2126 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00413 495 362 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00412 424 2115 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00411 424 2105 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00410 2044 2058 424 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00409 2044 424 620 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00408 2044 429 362 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00407 415 2126 418 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00406 2044 415 416 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00405 418 1464 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00404 2044 386 344 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00403 344 474 343 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00402 479 402 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00401 2044 399 402 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00400 350 348 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00399 402 1457 350 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00398 345 1899 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00397 2044 1764 345 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00396 2044 396 345 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00395 345 1457 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00394 394 1581 395 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00393 2044 394 396 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00392 395 911 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00391 2044 397 399 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00390 347 596 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00389 346 345 347 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00388 397 390 346 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00387 408 411 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00386 2044 2125 407 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00385 409 407 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 410 408 409 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00383 413 2125 410 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 2044 411 413 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 386 387 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 387 389 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00379 2044 1884 387 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00378 391 389 390 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00377 390 1898 391 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00376 391 1884 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00375 411 1464 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00374 2044 1884 411 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00373 2044 334 381 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00372 2044 576 389 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00371 2044 2055 382 2044 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00370 376 1764 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00369 383 410 336 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00368 336 2055 378 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00367 378 382 335 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00366 335 381 383 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00365 2044 1764 383 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00364 379 376 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00363 378 377 379 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00362 2044 378 1538 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00361 576 371 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00360 371 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00359 2044 2108 371 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00358 2044 1457 1757 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00357 2044 389 337 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00356 337 2115 453 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00355 330 332 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00354 2044 2058 332 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00353 264 1293 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00352 332 2108 264 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00351 2044 325 262 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00350 262 323 261 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00349 261 330 324 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00348 2044 2122 263 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00347 263 1293 355 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00346 325 326 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00345 326 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00344 2044 906 326 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00343 824 328 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00342 328 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00341 2044 355 328 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00340 319 322 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00339 322 720 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00338 2044 1753 322 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00337 254 507 316 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00336 316 313 254 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00335 254 1753 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 2044 906 255 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00333 255 1581 318 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00332 2044 411 312 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00331 313 312 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00330 2044 310 313 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00329 2044 1177 260 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00328 260 318 259 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00327 259 1884 320 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00326 2044 324 257 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00325 257 320 258 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00324 258 315 256 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00323 256 316 317 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00322 308 2122 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00321 2044 1899 308 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00320 306 304 253 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00319 2044 306 305 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00318 253 698 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00317 301 302 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00316 2044 319 302 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00315 252 1581 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00314 302 1884 252 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00313 2044 308 1018 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00312 2044 307 698 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00311 307 308 2044 2044 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00310 294 583 244 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00309 2044 294 304 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00308 244 1884 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00307 291 293 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00306 293 304 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00305 2044 1898 293 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00304 2044 343 246 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 246 295 247 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00302 247 297 245 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 245 301 298 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00300 2044 2058 249 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00299 249 296 248 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00298 248 423 297 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00297 251 317 299 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00296 2044 1849 251 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00295 250 1764 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00294 299 298 250 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00293 2044 299 348 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 2044 284 279 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 240 578 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 241 290 240 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 284 280 241 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00288 289 386 242 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00287 2044 289 287 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00286 242 1753 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00285 243 291 290 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00284 290 287 243 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00283 243 1764 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00282 286 281 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00281 2044 1457 286 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00280 2044 464 286 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00279 286 1899 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00278 2044 1849 1764 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 272 278 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 278 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00275 2044 2115 278 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00274 2044 272 273 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00273 2044 270 560 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00272 238 1753 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00271 239 272 238 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00270 270 266 239 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00269 2044 2108 236 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 236 2058 334 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 280 1541 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00266 2044 1757 280 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00265 2044 266 280 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00264 280 1899 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00263 265 334 237 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 2044 265 266 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 237 911 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 2044 310 227 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00259 227 720 1434 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00258 2044 230 1673 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00257 720 234 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00256 234 2126 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00255 2044 1189 234 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00254 229 2125 228 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00253 2044 229 230 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00252 228 2122 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00251 1189 232 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00250 232 2123 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00249 2044 1898 232 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00248 214 215 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00247 215 355 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00246 2044 2105 215 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00245 218 217 315 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 315 220 218 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 218 2058 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00242 212 2123 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00241 2044 2122 208 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00240 210 208 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00239 423 212 210 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00238 211 2122 423 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 2044 2123 211 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 2044 214 217 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00235 224 2113 223 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 2044 230 225 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00233 223 2058 226 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 225 2105 224 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 2044 226 221 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 2044 310 222 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 222 1673 220 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00228 220 2108 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00227 2044 205 203 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00226 206 203 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00225 2044 1189 206 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00224 2044 1581 207 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00223 207 2126 205 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00222 201 1018 202 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00221 202 205 201 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00220 2044 200 202 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00219 199 201 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 2044 206 200 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 198 195 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00216 2044 1673 198 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00215 177 2058 176 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00214 2044 177 281 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 176 198 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 192 390 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00211 2044 1899 192 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00210 192 1884 191 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00209 191 199 192 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00208 2044 191 477 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 2044 583 193 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 193 1899 296 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00205 583 196 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 196 195 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00203 2044 2126 196 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00202 190 1899 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00201 190 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00200 2044 198 190 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00199 2044 190 295 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 2044 2108 178 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 178 2126 179 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 2044 186 187 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00195 187 683 184 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00194 184 1884 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00193 2044 1581 185 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 185 1898 186 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00191 235 174 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00190 2044 279 174 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00189 175 182 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00188 174 1541 175 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00187 180 179 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00186 181 2113 683 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00185 2044 180 181 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00184 1068 164 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 2044 162 164 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00182 163 168 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00181 164 2058 163 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00180 2044 171 377 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 2044 167 166 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00178 166 273 2044 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00177 171 2055 172 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00176 172 169 2044 2044 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00175 166 1753 171 2044 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00174 161 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00173 2044 2113 160 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00172 159 160 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 168 161 159 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 158 2113 168 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 2044 2125 158 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 2044 168 173 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 2044 272 162 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 2044 2122 101 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00165 101 2055 152 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00164 2044 2122 1898 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00163 1898 2122 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 2044 2122 1898 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 1898 2122 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00160 2044 2108 99 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 99 2113 98 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 98 1189 148 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00157 155 720 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00156 2044 2105 155 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00155 323 195 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00154 2044 152 323 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00153 2044 150 1293 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 2044 2108 100 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 100 1899 363 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 102 2108 154 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 154 310 102 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00148 102 720 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 2044 363 149 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 146 149 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00145 146 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00144 2044 2055 146 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00143 2044 146 144 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 97 359 143 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 143 221 97 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 97 2055 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 2044 2113 96 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 96 362 141 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 133 1884 94 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00136 94 214 133 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00135 2044 137 94 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00134 134 133 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00133 2044 206 137 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00132 138 140 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00131 2044 144 140 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00130 95 141 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00129 140 2058 95 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00128 127 126 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00127 89 150 128 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 2044 127 89 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 2044 134 93 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 93 143 92 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00123 92 130 131 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00122 2044 129 91 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00121 91 128 90 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 90 138 130 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 129 1764 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00118 2044 122 129 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00117 150 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00116 2044 1899 150 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00115 121 1898 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00114 88 453 122 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 2044 121 88 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 2044 390 116 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 86 184 117 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 117 119 86 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 86 2055 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 114 179 85 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 85 2113 114 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00106 2044 116 85 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00105 113 114 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 120 122 87 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 2044 120 119 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 87 1884 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 82 2058 169 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 169 173 82 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 82 107 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00098 109 2058 83 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 2044 109 167 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 83 110 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 2044 107 81 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 81 126 443 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 112 2058 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00092 84 110 126 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 2044 112 84 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 104 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00089 2044 2113 103 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00088 79 103 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 110 104 79 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 80 2113 110 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 2044 2108 80 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00084 68 155 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00083 67 310 69 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 2044 68 67 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 2044 2055 1753 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 2044 2113 76 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 76 2058 75 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 75 155 74 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 310 70 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 70 2125 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00075 2044 1018 70 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00074 2044 310 73 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 73 77 72 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 72 74 71 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 78 1018 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00070 78 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 2044 2058 78 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00068 2044 78 77 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 2044 65 62 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 66 148 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 64 2058 66 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 65 69 64 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 2044 154 60 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00062 60 61 59 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00061 2044 61 63 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00060 59 63 58 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00059 58 69 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00058 57 59 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 61 56 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 56 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00055 2044 2058 56 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 53 71 54 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 2044 53 52 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 54 1753 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 50 305 51 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00050 51 62 50 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00049 2044 2055 51 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00048 49 50 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 1282 55 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 55 2113 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 2044 1884 55 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00044 2044 42 195 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 47 49 48 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 48 52 47 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 47 1764 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 2044 1189 46 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 46 2055 45 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 45 1282 43 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 43 42 44 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 2044 1457 35 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 35 131 34 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 40 44 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 39 272 41 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 2044 40 39 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 2044 48 32 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 32 36 33 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 33 31 30 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 30 34 182 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 2044 1849 38 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 38 57 37 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 37 41 36 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 22 2058 21 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 2044 22 23 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 21 1898 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 2044 1849 28 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 28 117 26 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 26 24 27 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 2044 286 29 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 29 27 31 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 25 23 24 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 24 113 25 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 25 1753 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 2044 2058 1884 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 14 1884 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 13 18 107 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 2044 14 13 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 42 20 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 20 2108 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 2044 2113 20 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 17 42 2044 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 2044 2125 16 2044 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 15 16 2044 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 18 17 15 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 19 2125 18 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 2044 42 19 2044 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C2146 1 2044 9.7e-15
C2132 14 2044 1.662e-14
C2130 16 2044 2.596e-14
C2129 17 2044 2.16e-14
C2128 18 2044 6.06e-14
C2126 20 2044 1.8635e-14
C2124 22 2044 1.8635e-14
C2123 23 2044 5.203e-14
C2122 24 2044 5.192e-14
C2121 25 2044 4.11e-15
C2119 27 2044 5.75e-14
C2115 31 2044 5.406e-14
C2112 34 2044 5.586e-14
C2110 36 2044 6.09e-14
C2106 40 2044 1.662e-14
C2105 41 2044 6.186e-14
C2104 42 2044 1.8464e-13
C2102 44 2044 6.325e-14
C2099 47 2044 4.11e-15
C2098 48 2044 8.912e-14
C2097 49 2044 4.727e-14
C2096 50 2044 1.853e-14
C2095 51 2044 4.11e-15
C2094 52 2044 5.593e-14
C2093 53 2044 1.8635e-14
C2091 55 2044 1.8635e-14
C2090 56 2044 1.8635e-14
C2089 57 2044 1.3824e-13
C2087 59 2044 1.932e-14
C2085 61 2044 7.196e-14
C2084 62 2044 9.121e-14
C2083 63 2044 2.356e-14
C2081 65 2044 2.605e-14
C2078 68 2044 1.662e-14
C2077 69 2044 8.813e-14
C2076 70 2044 1.8635e-14
C2075 71 2044 1.1771e-13
C2072 74 2044 5.76e-14
C2069 77 2044 6.912e-14
C2068 78 2044 2.455e-14
C2064 82 2044 4.11e-15
C2061 85 2044 4.11e-15
C2060 86 2044 4.11e-15
C2052 94 2044 4.11e-15
C2049 97 2044 4.11e-15
C2044 102 2044 4.11e-15
C2042 103 2044 2.596e-14
C2041 104 2044 2.16e-14
C2040 105 2044 9.7e-15
C2039 106 2044 6.05e-15
C2038 107 2044 1.029e-13
C2036 109 2044 1.8635e-14
C2035 110 2044 1.0597e-13
C2034 111 2044 6.05e-15
C2033 112 2044 1.662e-14
C2032 113 2044 5.477e-14
C2031 114 2044 1.853e-14
C2029 116 2044 5.525e-14
C2028 117 2044 6.612e-14
C2026 119 2044 4.633e-14
C2025 120 2044 1.8635e-14
C2024 121 2044 1.662e-14
C2023 122 2044 7.323e-14
C2019 126 2044 1.6381e-13
C2018 127 2044 1.662e-14
C2017 128 2044 5.686e-14
C2016 129 2044 6.591e-14
C2015 130 2044 5.76e-14
C2014 131 2044 9.278e-14
C2012 133 2044 1.853e-14
C2011 134 2044 6.307e-14
C2008 137 2044 5.525e-14
C2007 138 2044 8.612e-14
C2006 139 2044 6.05e-15
C2005 140 2044 1.767e-14
C2004 141 2044 4.731e-14
C2002 143 2044 9.372e-14
C2001 144 2044 7.633e-14
C1999 146 2044 2.455e-14
C1997 148 2044 5.703e-14
C1996 149 2044 5.259e-14
C1995 150 2044 2.0153e-13
C1993 152 2044 5.016e-14
C1991 154 2044 1.1581e-13
C1990 155 2044 1.2717e-13
C1988 157 2044 9.7e-15
C1985 160 2044 2.596e-14
C1984 161 2044 2.16e-14
C1983 162 2044 5.285e-14
C1981 164 2044 1.767e-14
C1979 166 2044 4.11e-15
C1978 167 2044 5.218e-14
C1977 168 2044 9.346e-14
C1976 169 2044 5.372e-14
C1975 170 2044 8.58e-15
C1974 171 2044 2.299e-14
C1972 173 2044 5.529e-14
C1971 174 2044 1.767e-14
C1968 177 2044 1.8635e-14
C1966 179 2044 8.256e-14
C1965 180 2044 1.662e-14
C1963 182 2044 9.761e-14
C1962 183 2044 6.05e-15
C1961 184 2044 5.005e-14
C1959 186 2044 4.341e-14
C1955 190 2044 2.455e-14
C1954 191 2044 2.639e-14
C1953 192 2044 7.43e-15
C1950 195 2044 2.3621e-13
C1949 196 2044 1.8635e-14
C1947 198 2044 1.471e-13
C1946 199 2044 7.427e-14
C1945 200 2044 5.525e-14
C1944 201 2044 1.853e-14
C1943 202 2044 4.11e-15
C1942 203 2044 1.677e-14
C1940 205 2044 9.292e-14
C1939 206 2044 8.544e-14
C1937 208 2044 2.596e-14
C1936 209 2044 9.7e-15
C1933 212 2044 2.16e-14
C1931 214 2044 1.2168e-13
C1930 215 2044 1.8635e-14
C1928 217 2044 5.019e-14
C1927 218 2044 4.11e-15
C1926 219 2044 6.05e-15
C1925 220 2044 4.747e-14
C1924 221 2044 9.273e-14
C1919 226 2044 2.306e-14
C1916 229 2044 1.8635e-14
C1915 230 2044 8.269e-14
C1913 232 2044 1.8635e-14
C1910 234 2044 1.8635e-14
C1909 235 2044 7.247e-14
C1901 243 2044 4.11e-15
C1890 254 2044 4.11e-15
C1878 265 2044 1.8635e-14
C1877 266 2044 8.161e-14
C1873 270 2044 2.605e-14
C1871 272 2044 2.4557e-13
C1870 273 2044 4.326e-14
C1867 276 2044 7.56e-15
C1865 278 2044 1.8635e-14
C1864 279 2044 6.101e-14
C1863 280 2044 6.751e-14
C1862 281 2044 5.188e-14
C1859 284 2044 2.605e-14
C1857 286 2044 9.909e-14
C1856 287 2044 5.641e-14
C1854 289 2044 1.8635e-14
C1853 290 2044 5.957e-14
C1852 291 2044 4.391e-14
C1850 293 2044 1.8635e-14
C1849 294 2044 1.8635e-14
C1848 295 2044 6.782e-14
C1847 296 2044 5.686e-14
C1846 297 2044 5.58e-14
C1845 298 2044 6.911e-14
C1844 299 2044 2.445e-14
C1843 300 2044 7.43e-15
C1842 301 2044 7.892e-14
C1841 302 2044 1.767e-14
C1840 303 2044 6.05e-15
C1839 304 2044 1.3252e-13
C1838 305 2044 8.281e-14
C1837 306 2044 1.8635e-14
C1836 307 2044 1.568e-14
C1835 308 2044 8.616e-14
C1833 310 2044 3.0198e-13
C1831 312 2044 1.677e-14
C1830 313 2044 5.539e-14
C1828 315 2044 5.204e-14
C1827 316 2044 6.032e-14
C1826 317 2044 1.1591e-13
C1825 318 2044 7.294e-14
C1824 319 2044 1.2817e-13
C1823 320 2044 5.37e-14
C1821 322 2044 1.8635e-14
C1820 323 2044 6.788e-14
C1819 324 2044 6.84e-14
C1818 325 2044 5.251e-14
C1817 326 2044 1.8635e-14
C1815 328 2044 1.8635e-14
C1813 330 2044 7.892e-14
C1812 331 2044 6.05e-15
C1811 332 2044 1.767e-14
C1809 334 2044 8.168e-14
C1800 343 2044 5.826e-14
C1798 345 2044 6.121e-14
C1795 348 2044 5.233e-14
C1794 349 2044 6.05e-15
C1792 351 2044 9.7e-15
C1788 355 2044 2.0981e-13
C1784 359 2044 7.531e-14
C1781 362 2044 1.332e-13
C1780 363 2044 1.0955e-13
C1775 368 2044 5.525e-14
C1774 369 2044 4.11e-15
C1771 371 2044 1.8635e-14
C1769 373 2044 7.56e-15
C1766 376 2044 2.378e-14
C1765 377 2044 6.722e-14
C1764 378 2044 3.608e-14
C1761 381 2044 5.808e-14
C1760 382 2044 2.128e-14
C1759 383 2044 7.56e-15
C1756 386 2044 1.144e-13
C1755 387 2044 1.8635e-14
C1753 389 2044 1.1949e-13
C1752 390 2044 1.8557e-13
C1751 391 2044 4.11e-15
C1748 394 2044 1.8635e-14
C1746 396 2044 5.278e-14
C1745 397 2044 2.605e-14
C1744 398 2044 4.11e-15
C1743 399 2044 6.221e-14
C1740 402 2044 1.767e-14
C1737 405 2044 7.56e-15
C1735 407 2044 2.596e-14
C1734 408 2044 2.16e-14
C1732 410 2044 1.3862e-13
C1731 411 2044 1.2962e-13
C1727 415 2044 1.8635e-14
C1726 416 2044 5.203e-14
C1725 417 2044 4.11e-15
C1723 419 2044 2.455e-14
C1719 423 2044 1.7315e-13
C1718 424 2044 2.455e-14
C1716 426 2044 4.11e-15
C1713 429 2044 1.0089e-13
C1709 433 2044 6.82e-14
C1708 434 2044 5.63e-14
C1705 437 2044 1.853e-14
C1704 438 2044 5.492e-14
C1702 440 2044 4.11e-15
C1698 443 2044 1.046e-13
C1697 444 2044 2.378e-14
C1695 446 2044 2.128e-14
C1694 447 2044 3.608e-14
C1692 449 2044 7.56e-15
C1690 451 2044 2.596e-14
C1689 452 2044 5.654e-14
C1688 453 2044 1.8257e-13
C1687 454 2044 9.7e-15
C1686 455 2044 2.16e-14
C1685 456 2044 1.8635e-14
C1684 457 2044 8.289e-14
C1681 460 2044 1.677e-14
C1680 461 2044 5.581e-14
C1677 464 2044 6.862e-14
C1676 465 2044 8.745e-14
C1675 466 2044 1.8635e-14
C1674 467 2044 1.662e-14
C1673 468 2044 5.255e-14
C1672 469 2044 5.436e-14
C1670 471 2044 2.455e-14
C1667 474 2044 8.437e-14
C1665 476 2044 5.292e-14
C1664 477 2044 8.176e-14
C1662 479 2044 5.71e-14
C1661 480 2044 1.3221e-13
C1659 482 2044 2.378e-14
C1658 483 2044 2.128e-14
C1656 485 2044 3.608e-14
C1654 487 2044 7.56e-15
C1653 488 2044 4.424e-14
C1652 489 2044 2.445e-14
C1651 490 2044 7.43e-15
C1650 491 2044 1.0729e-13
C1648 493 2044 1.853e-14
C1647 494 2044 5.953e-14
C1646 495 2044 7.462e-14
C1644 497 2044 1.0003e-13
C1643 498 2044 4.921e-14
C1642 499 2044 1.767e-14
C1641 500 2044 6.05e-15
C1640 501 2044 7.292e-14
C1639 502 2044 1.1969e-13
C1638 503 2044 7.335e-14
C1636 505 2044 1.8635e-14
C1634 507 2044 6.667e-14
C1631 510 2044 8.58e-15
C1630 511 2044 5.725e-14
C1629 512 2044 1.1703e-13
C1627 514 2044 1.677e-14
C1626 515 2044 6.223e-14
C1625 516 2044 6.586e-14
C1623 518 2044 7.649e-14
C1622 519 2044 1.2916e-13
C1620 521 2044 1.8635e-14
C1619 522 2044 5.231e-14
C1618 523 2044 6.05e-15
C1617 524 2044 4.987e-14
C1616 525 2044 1.386e-13
C1614 527 2044 1.7683e-13
C1613 528 2044 2.605e-14
C1612 529 2044 4.755e-14
C1611 530 2044 9.7e-15
C1607 534 2044 6.05e-15
C1604 537 2044 8.58e-15
C1602 539 2044 6.05e-15
C1596 545 2044 6.05e-15
C1595 546 2044 7.43e-15
C1592 549 2044 6.05e-15
C1591 550 2044 6.05e-15
C1587 554 2044 6.05e-15
C1583 557 2044 2.596e-14
C1580 560 2044 7.995e-14
C1579 561 2044 2.16e-14
C1577 563 2044 5.839e-14
C1575 565 2044 2.72e-14
C1574 566 2044 5.103e-14
C1573 567 2044 1.1999e-13
C1571 569 2044 4.11e-15
C1570 570 2044 7.43e-15
C1569 571 2044 4.11e-15
C1568 572 2044 1.853e-14
C1566 574 2044 4.415e-14
C1564 576 2044 1.8929e-13
C1563 577 2044 4.11e-15
C1562 578 2044 8.555e-14
C1561 579 2044 4.352e-14
C1560 580 2044 5.957e-14
C1558 582 2044 1.767e-14
C1557 583 2044 1.8249e-13
C1556 584 2044 4.11e-15
C1555 585 2044 1.853e-14
C1552 588 2044 8.863e-14
C1551 589 2044 8.977e-14
C1550 590 2044 5.026e-14
C1548 592 2044 1.8635e-14
C1545 595 2044 1.767e-14
C1544 596 2044 7.835e-14
C1543 597 2044 4.11e-15
C1542 598 2044 8.236e-14
C1540 600 2044 6.135e-14
C1538 602 2044 5.175e-14
C1537 603 2044 2.445e-14
C1529 611 2044 2.306e-14
C1528 612 2044 1.6463e-13
C1522 618 2044 8.467e-14
C1520 620 2044 1.2621e-13
C1519 621 2044 6.911e-14
C1517 623 2044 7.236e-14
C1516 624 2044 4.11e-15
C1514 626 2044 1.8635e-14
C1512 628 2044 5.477e-14
C1511 629 2044 1.767e-14
C1506 634 2044 1.2163e-13
C1504 636 2044 1.8635e-14
C1502 638 2044 5.201e-14
C1499 641 2044 2.605e-14
C1498 642 2044 5.001e-14
C1491 649 2044 8.387e-14
C1490 650 2044 8.337e-14
C1489 651 2044 9.032e-14
C1488 652 2044 4.11e-15
C1484 656 2044 4.477e-14
C1481 659 2044 5.601e-14
C1479 661 2044 1.8635e-14
C1476 663 2044 1.2147e-13
C1475 664 2044 5.94e-14
C1474 665 2044 1.662e-14
C1473 666 2044 1.8635e-14
C1472 667 2044 7.809e-14
C1471 668 2044 5.893e-14
C1469 670 2044 2.639e-14
C1467 672 2044 1.8635e-14
C1465 674 2044 4.987e-14
C1464 675 2044 6.05e-15
C1463 676 2044 1.767e-14
C1462 677 2044 5.312e-14
C1461 678 2044 1.8635e-14
C1458 681 2044 1.1905e-13
C1457 682 2044 1.8635e-14
C1456 683 2044 1.3305e-13
C1455 684 2044 5.876e-14
C1453 686 2044 5.781e-14
C1451 688 2044 6.05e-15
C1450 689 2044 4.747e-14
C1449 690 2044 6.332e-14
C1448 691 2044 9.09e-14
C1447 692 2044 5.728e-14
C1446 693 2044 6.071e-14
C1445 694 2044 7.43e-15
C1444 695 2044 2.445e-14
C1443 696 2044 1.8635e-14
C1442 697 2044 5.358e-14
C1441 698 2044 1.2488e-13
C1440 699 2044 1.662e-14
C1439 700 2044 2.605e-14
C1438 701 2044 5.243e-14
C1437 702 2044 9.72e-14
C1436 703 2044 1.8635e-14
C1434 705 2044 6.186e-14
C1433 706 2044 1.8635e-14
C1431 708 2044 5.396e-14
C1430 709 2044 5.62e-14
C1429 710 2044 6.427e-14
C1426 713 2044 2.455e-14
C1424 715 2044 1.3918e-13
C1423 716 2044 1.0078e-13
C1422 717 2044 5.337e-14
C1421 718 2044 2.306e-14
C1420 719 2044 5.256e-14
C1419 720 2044 3.3992e-13
C1417 722 2044 6.05e-15
C1410 729 2044 9.37e-15
C1409 730 2044 7.33e-15
C1408 731 2044 1.154e-14
C1407 732 2044 6.05e-15
C1400 739 2044 9.96e-15
C1398 741 2044 6.05e-15
C1396 743 2044 7.43e-15
C1393 745 2044 1.8635e-14
C1391 747 2044 1.8635e-14
C1389 749 2044 4.11e-15
C1388 750 2044 9.21e-14
C1387 751 2044 5.473e-14
C1386 752 2044 6.467e-14
C1385 753 2044 4.11e-15
C1384 754 2044 4.179e-14
C1383 755 2044 6.501e-14
C1382 756 2044 7.352e-14
C1380 758 2044 1.8635e-14
C1379 759 2044 4.926e-14
C1377 761 2044 7.127e-14
C1376 762 2044 4.11e-15
C1372 766 2044 1.9199e-13
C1369 769 2044 2.605e-14
C1368 770 2044 5.745e-14
C1367 771 2044 8.63e-14
C1366 772 2044 4.11e-15
C1365 773 2044 9.708e-14
C1362 776 2044 1.8635e-14
C1358 780 2044 1.9813e-13
C1357 781 2044 4.11e-15
C1356 782 2044 8.784e-14
C1355 783 2044 4.11e-15
C1353 785 2044 5.291e-14
C1351 787 2044 6.908e-14
C1350 788 2044 5.102e-14
C1346 792 2044 3.405e-14
C1344 794 2044 6.047e-14
C1343 795 2044 1.767e-14
C1339 799 2044 5.772e-14
C1338 800 2044 4.11e-15
C1336 802 2044 1.2348e-13
C1335 803 2044 1.8635e-14
C1334 804 2044 7.43e-15
C1333 805 2044 4.907e-14
C1332 806 2044 6.525e-14
C1331 807 2044 8.823e-14
C1330 808 2044 4.11e-15
C1329 809 2044 2.259e-14
C1324 814 2044 5.04e-14
C1320 818 2044 5.346e-14
C1319 819 2044 1.8635e-14
C1318 820 2044 1.3835e-13
C1317 821 2044 4.11e-15
C1314 824 2044 1.0027e-13
C1312 826 2044 1.767e-14
C1311 827 2044 7.56e-15
C1308 830 2044 4.541e-14
C1307 831 2044 1.8635e-14
C1304 834 2044 5.529e-14
C1303 835 2044 9.658e-14
C1302 836 2044 2.445e-14
C1295 843 2044 2.6525e-13
C1292 846 2044 6.48e-14
C1291 847 2044 6.872e-14
C1290 848 2044 1.0028e-13
C1289 849 2044 5.654e-14
C1288 850 2044 5.94e-14
C1286 852 2044 7.43e-15
C1284 854 2044 6.44e-14
C1283 855 2044 6.05e-15
C1282 856 2044 2.9509e-13
C1280 858 2044 4.731e-14
C1279 859 2044 1.7144e-13
C1276 862 2044 6.286e-14
C1274 864 2044 2.356e-14
C1270 867 2044 2.455e-14
C1267 870 2044 5.747e-14
C1266 871 2044 1.0179e-13
C1264 873 2044 1.677e-14
C1263 874 2044 8.101e-14
C1261 876 2044 7.76e-15
C1260 877 2044 9.7e-15
C1258 879 2044 6.209e-14
C1257 880 2044 4.771e-14
C1255 882 2044 1.8635e-14
C1254 883 2044 9.7e-15
C1252 885 2044 5.516e-14
C1250 887 2044 8.58e-15
C1249 888 2044 1.8635e-14
C1248 889 2044 8.674e-14
C1245 892 2044 2.445e-14
C1244 893 2044 6.732e-14
C1242 895 2044 7.56e-15
C1241 896 2044 1.8635e-14
C1240 897 2044 5.396e-14
C1236 901 2044 5.853e-14
C1235 902 2044 1.767e-14
C1232 905 2044 1.8635e-14
C1231 906 2044 2.2792e-13
C1228 909 2044 1.932e-14
C1227 910 2044 6.05e-15
C1226 911 2044 5.5014e-13
C1223 914 2044 8.326e-14
C1220 917 2044 2.378e-14
C1219 918 2044 6.096e-14
C1218 919 2044 2.128e-14
C1216 921 2044 3.608e-14
C1215 922 2044 7.56e-15
C1212 925 2044 2.16e-14
C1211 926 2044 1.2812e-13
C1210 927 2044 2.596e-14
C1209 928 2044 7.76e-15
C1207 930 2044 7.56e-15
C1204 932 2044 2.596e-14
C1203 933 2044 7.43e-15
C1201 935 2044 5.049e-14
C1199 937 2044 2.16e-14
C1197 939 2044 9.459e-14
C1196 940 2044 7.86e-14
C1194 942 2044 1.8635e-14
C1192 944 2044 2.596e-14
C1190 946 2044 2.16e-14
C1189 947 2044 1.1397e-13
C1188 948 2044 1.8635e-14
C1186 950 2044 2.596e-14
C1185 951 2044 1.1931e-13
C1183 953 2044 2.16e-14
C1180 956 2044 5.1e-14
C1178 958 2044 1.662e-14
C1176 960 2044 1.8635e-14
C1175 961 2044 6.972e-14
C1174 962 2044 5.248e-14
C1172 964 2044 2.299e-14
C1171 965 2044 4.11e-15
C1167 969 2044 2.605e-14
C1166 970 2044 5.178e-14
C1165 971 2044 1.0456e-13
C1162 974 2044 8.64e-14
C1161 975 2044 1.0794e-13
C1159 977 2044 2.378e-14
C1157 979 2044 7.424e-14
C1156 980 2044 3.608e-14
C1154 982 2044 7.56e-15
C1153 983 2044 2.128e-14
C1152 984 2044 1.5263e-13
C1150 986 2044 1.8635e-14
C1149 987 2044 8.014e-14
C1147 989 2044 1.8234e-13
C1146 990 2044 1.8635e-14
C1145 991 2044 1.662e-14
C1143 993 2044 1.3662e-13
C1141 995 2044 1.8635e-14
C1140 996 2044 7.176e-14
C1139 997 2044 2.3186e-13
C1138 998 2044 1.8635e-14
C1136 1000 2044 1.767e-14
C1135 1001 2044 1.8635e-14
C1133 1003 2044 1.677e-14
C1132 1004 2044 9.829e-14
C1131 1005 2044 1.0069e-13
C1130 1006 2044 2.2199e-13
C1129 1007 2044 1.662e-14
C1127 1009 2044 6.344e-14
C1126 1010 2044 7.052e-14
C1124 1012 2044 2.378e-14
C1122 1014 2044 7.56e-15
C1121 1015 2044 3.608e-14
C1119 1017 2044 2.128e-14
C1118 1018 2044 5.0528e-13
C1117 1019 2044 1.8635e-14
C1111 1025 2044 7.56e-15
C1105 1031 2044 7.56e-15
C1100 1036 2044 7.56e-15
C1094 1042 2044 7.56e-15
C1091 1045 2044 4.11e-15
C1088 1048 2044 4.11e-15
C1085 1051 2044 4.11e-15
C1084 1052 2044 4.11e-15
C1080 1056 2044 4.11e-15
C1076 1059 2044 9.7e-15
C1075 1060 2044 2.596e-14
C1073 1062 2044 2.16e-14
C1070 1065 2044 7.56e-15
C1069 1066 2044 2.128e-14
C1068 1067 2044 2.378e-14
C1067 1068 2044 1.7134e-13
C1066 1069 2044 4.958e-14
C1063 1072 2044 3.608e-14
C1061 1074 2044 2.596e-14
C1060 1075 2044 7.56e-15
C1057 1078 2044 9.618e-14
C1056 1079 2044 2.16e-14
C1055 1080 2044 7.76e-15
C1054 1081 2044 8.151e-14
C1053 1082 2044 1.1026e-13
C1052 1083 2044 1.8635e-14
C1049 1086 2044 2.128e-14
C1048 1087 2044 2.378e-14
C1046 1089 2044 3.608e-14
C1043 1092 2044 7.76e-15
C1042 1093 2044 7.56e-15
C1041 1094 2044 3.864e-14
C1039 1096 2044 9.515e-14
C1038 1097 2044 1.8635e-14
C1036 1099 2044 8.494e-14
C1035 1100 2044 1.662e-14
C1034 1101 2044 1.8635e-14
C1030 1105 2044 2.128e-14
C1029 1106 2044 2.378e-14
C1028 1107 2044 6.082e-14
C1026 1109 2044 7.56e-15
C1025 1110 2044 3.608e-14
C1022 1113 2044 5.686e-14
C1019 1116 2044 7.56e-15
C1017 1118 2044 6.221e-14
C1016 1119 2044 8.29e-14
C1015 1120 2044 2.0013e-13
C1014 1121 2044 1.767e-14
C1013 1122 2044 6.05e-15
C1010 1125 2044 7.56e-15
C1009 1126 2044 2.128e-14
C1008 1127 2044 2.378e-14
C1007 1128 2044 7.34e-14
C1005 1130 2044 3.608e-14
C1002 1133 2044 7.56e-15
C998 1137 2044 7.56e-15
C997 1138 2044 1.513e-13
C996 1139 2044 1.8635e-14
C995 1140 2044 1.853e-14
C993 1142 2044 1.7058e-13
C992 1143 2044 5.113e-14
C990 1145 2044 5.057e-14
C987 1148 2044 7.56e-15
C985 1150 2044 5.601e-14
C984 1151 2044 2.605e-14
C983 1152 2044 4.95e-14
C982 1153 2044 6.302e-14
C981 1154 2044 2.299e-14
C977 1158 2044 8.58e-15
C975 1160 2044 1.8635e-14
C973 1162 2044 7.379e-14
C971 1164 2044 3.5573e-13
C970 1165 2044 2.299e-14
C967 1168 2044 1.5034e-13
C966 1169 2044 8.58e-15
C965 1170 2044 1.7014e-13
C962 1173 2044 6.05e-15
C961 1174 2044 1.767e-14
C960 1175 2044 4.767e-14
C959 1176 2044 6.05e-15
C958 1177 2044 2.0848e-13
C957 1178 2044 1.767e-14
C956 1179 2044 5.117e-14
C955 1180 2044 6.05e-15
C952 1183 2044 1.0388e-13
C951 1184 2044 5.773e-14
C948 1187 2044 8.529e-14
C947 1188 2044 8.58e-15
C946 1189 2044 5.5193e-13
C945 1190 2044 8.003e-14
C944 1191 2044 1.767e-14
C943 1192 2044 6.05e-15
C941 1193 2044 6.05e-15
C940 1194 2044 2.757e-14
C938 1196 2044 2.378e-14
C937 1197 2044 4.506e-14
C936 1198 2044 1.2802e-13
C935 1199 2044 3.608e-14
C933 1201 2044 7.56e-15
C932 1202 2044 2.128e-14
C930 1204 2044 2.9396e-13
C929 1205 2044 5.065e-14
C928 1206 2044 4.11e-15
C927 1207 2044 1.853e-14
C926 1208 2044 1.8635e-14
C925 1209 2044 1.4034e-13
C923 1211 2044 1.2114e-13
C921 1213 2044 6.282e-14
C920 1214 2044 1.0211e-13
C919 1215 2044 1.853e-14
C918 1216 2044 4.11e-15
C917 1217 2044 2.596e-14
C915 1219 2044 2.16e-14
C913 1221 2044 4.993e-14
C912 1222 2044 5.717e-14
C911 1223 2044 1.853e-14
C910 1224 2044 4.11e-15
C909 1225 2044 5.057e-14
C908 1226 2044 6.28e-14
C906 1228 2044 5.327e-14
C905 1229 2044 2.356e-14
C903 1231 2044 1.932e-14
C901 1233 2044 6.452e-14
C899 1235 2044 5.684e-14
C898 1236 2044 1.1632e-13
C897 1237 2044 2.378e-14
C895 1239 2044 2.128e-14
C894 1240 2044 7.56e-15
C893 1241 2044 3.608e-14
C891 1243 2044 1.7373e-13
C889 1245 2044 2.378e-14
C888 1246 2044 6.81e-14
C887 1247 2044 3.608e-14
C885 1249 2044 2.128e-14
C883 1251 2044 7.56e-15
C882 1252 2044 5.122e-14
C880 1254 2044 1.573e-13
C879 1255 2044 2.378e-14
C878 1256 2044 7.56e-15
C875 1259 2044 3.608e-14
C874 1260 2044 2.128e-14
C873 1261 2044 5.466e-14
C871 1263 2044 1.244e-13
C870 1264 2044 2.378e-14
C868 1266 2044 7.56e-15
C867 1267 2044 3.608e-14
C865 1269 2044 2.128e-14
C864 1270 2044 3.992e-14
C863 1271 2044 4.11e-15
C862 1272 2044 1.853e-14
C861 1273 2044 2.1565e-13
C860 1274 2044 4.11e-15
C859 1275 2044 5.447e-14
C858 1276 2044 1.0076e-13
C857 1277 2044 4.11e-15
C855 1279 2044 4.611e-14
C854 1280 2044 2.5108e-13
C853 1281 2044 7.159e-14
C852 1282 2044 3.5218e-13
C851 1283 2044 7.43e-15
C850 1284 2044 6.013e-14
C849 1285 2044 1.767e-14
C847 1287 2044 5.405e-14
C846 1288 2044 5.057e-14
C845 1289 2044 4.11e-15
C844 1290 2044 1.0572e-13
C843 1291 2044 6.485e-14
C841 1293 2044 4.1687e-13
C840 1294 2044 5.211e-14
C839 1295 2044 1.767e-14
C835 1299 2044 7.56e-15
C831 1303 2044 4.11e-15
C825 1309 2044 4.11e-15
C824 1310 2044 4.11e-15
C820 1314 2044 7.56e-15
C819 1315 2044 4.11e-15
C815 1319 2044 7.56e-15
C810 1324 2044 7.56e-15
C803 1331 2044 7.56e-15
C802 1332 2044 4.11e-15
C795 1338 2044 2.378e-14
C794 1339 2044 5.9e-14
C792 1341 2044 2.128e-14
C790 1343 2044 3.608e-14
C788 1345 2044 7.56e-15
C787 1346 2044 2.2699e-13
C786 1347 2044 1.767e-14
C785 1348 2044 6.05e-15
C784 1349 2044 4.172e-14
C783 1350 2044 6.53e-14
C782 1351 2044 5.405e-14
C781 1352 2044 2.299e-14
C779 1354 2044 8.58e-15
C778 1355 2044 4.284e-14
C777 1356 2044 1.767e-14
C776 1357 2044 6.05e-15
C775 1358 2044 8.148e-14
C774 1359 2044 1.0929e-13
C773 1360 2044 5.405e-14
C772 1361 2044 1.767e-14
C771 1362 2044 6.05e-15
C770 1363 2044 6.418e-14
C769 1364 2044 1.8635e-14
C768 1365 2044 8.313e-14
C767 1366 2044 1.662e-14
C765 1368 2044 1.8635e-14
C760 1373 2044 1.5782e-13
C758 1375 2044 1.8635e-14
C757 1376 2044 7.56e-15
C755 1378 2044 5.554e-14
C751 1382 2044 2.128e-14
C750 1383 2044 2.378e-14
C749 1384 2044 5e-14
C747 1386 2044 3.608e-14
C746 1387 2044 7.56e-15
C744 1389 2044 7.56e-15
C742 1391 2044 1.2708e-13
C740 1393 2044 5.36e-14
C739 1394 2044 7.868e-14
C738 1395 2044 1.0908e-13
C737 1396 2044 2.128e-14
C736 1397 2044 2.378e-14
C735 1398 2044 1.0402e-13
C732 1401 2044 5.826e-14
C731 1402 2044 3.608e-14
C730 1403 2044 7.56e-15
C727 1406 2044 1.0198e-13
C726 1407 2044 5.769e-14
C722 1411 2044 7.56e-15
C721 1412 2044 2.128e-14
C720 1413 2044 2.378e-14
C718 1415 2044 3.608e-14
C716 1417 2044 4.642e-14
C715 1418 2044 7.56e-15
C714 1419 2044 3.9159e-13
C713 1420 2044 1.261e-13
C711 1422 2044 2.128e-14
C710 1423 2044 2.378e-14
C709 1424 2044 6.352e-14
C706 1427 2044 3.608e-14
C705 1428 2044 1.3703e-13
C704 1429 2044 3.864e-14
C703 1430 2044 7.56e-15
C702 1431 2044 1.4428e-13
C700 1433 2044 1.853e-14
C699 1434 2044 1.9452e-13
C698 1435 2044 4.453e-14
C695 1438 2044 2.7285e-14
C694 1439 2044 1.0992e-13
C693 1440 2044 7.076e-14
C692 1441 2044 5.567e-14
C689 1444 2044 1.932e-14
C688 1445 2044 2.356e-14
C687 1446 2044 7.467e-14
C683 1450 2044 4.11e-15
C681 1452 2044 4.11e-15
C680 1453 2044 7.101e-14
C678 1455 2044 4.11e-15
C677 1456 2044 5.733e-14
C676 1457 2044 7.789e-13
C674 1459 2044 4.11e-15
C673 1460 2044 6.933e-14
C671 1462 2044 4.11e-15
C670 1463 2044 4.637e-14
C669 1464 2044 3.8985e-13
C667 1466 2044 4.11e-15
C666 1467 2044 6.05e-15
C664 1469 2044 5.123e-14
C663 1470 2044 1.5975e-13
C660 1473 2044 7.662e-14
C659 1474 2044 5.645e-14
C658 1475 2044 6.05e-15
C656 1477 2044 5.803e-14
C654 1479 2044 6.06e-14
C652 1481 2044 2.378e-14
C651 1482 2044 3.608e-14
C649 1484 2044 2.128e-14
C648 1485 2044 7.56e-15
C646 1487 2044 7.412e-14
C645 1488 2044 6.98e-14
C643 1490 2044 2.378e-14
C641 1492 2044 1.212e-13
C640 1493 2044 7.56e-15
C639 1494 2044 2.128e-14
C637 1496 2044 3.608e-14
C635 1498 2044 4.11e-15
C634 1499 2044 6.128e-14
C632 1501 2044 4.11e-15
C631 1502 2044 6.05e-15
C629 1504 2044 6.754e-14
C628 1505 2044 8.42e-14
C626 1507 2044 2.378e-14
C625 1508 2044 5.002e-14
C622 1511 2044 3.608e-14
C621 1512 2044 7.56e-15
C620 1513 2044 2.128e-14
C618 1515 2044 4.266e-14
C616 1517 2044 1.574e-13
C615 1518 2044 4.11e-15
C613 1520 2044 4.11e-15
C612 1521 2044 1.677e-14
C611 1522 2044 1.1679e-13
C609 1524 2044 6.883e-14
C608 1525 2044 6.05e-15
C606 1527 2044 1.2985e-13
C604 1529 2044 5.617e-14
C601 1532 2044 1.4687e-13
C600 1533 2044 8.735e-14
C596 1536 2044 4.11e-15
C595 1537 2044 4.569e-14
C594 1538 2044 1.7061e-13
C593 1539 2044 5.892e-14
C592 1540 2044 5.072e-14
C591 1541 2044 6.25219e-13
C590 1542 2044 5.927e-14
C589 1543 2044 4.11e-15
C588 1544 2044 1.6228e-13
C587 1545 2044 1.853e-14
C586 1546 2044 6.575e-14
C585 1547 2044 4.11e-15
C584 1548 2044 1.853e-14
C583 1549 2044 4.11e-15
C582 1550 2044 1.853e-14
C581 1551 2044 1.853e-14
C579 1553 2044 2.3352e-13
C577 1555 2044 1.8635e-14
C573 1559 2044 7.56e-15
C572 1560 2044 1.8635e-14
C571 1561 2044 1.767e-14
C570 1562 2044 4.11e-15
C567 1565 2044 4.11e-15
C565 1567 2044 1.6056e-13
C563 1569 2044 1.1145e-13
C562 1570 2044 8.898e-14
C561 1571 2044 4.11e-15
C560 1572 2044 1.767e-14
C559 1573 2044 4.11e-15
C556 1576 2044 4.11e-15
C555 1577 2044 1.2693e-13
C554 1578 2044 4.11e-15
C553 1579 2044 6.759e-14
C551 1581 2044 6.3291e-13
C548 1584 2044 7.56e-15
C547 1585 2044 1.767e-14
C546 1586 2044 1.8635e-14
C544 1588 2044 4.11e-15
C543 1589 2044 1.8635e-14
C541 1591 2044 4.11e-15
C540 1592 2044 1.853e-14
C535 1596 2044 5.057e-14
C533 1598 2044 1.853e-14
C532 1599 2044 5.597e-14
C531 1600 2044 5.597e-14
C530 1601 2044 1.853e-14
C528 1603 2044 5.733e-14
C526 1605 2044 1.853e-14
C524 1607 2044 6.121e-14
C523 1608 2044 5.814e-14
C522 1609 2044 2.8006e-13
C521 1610 2044 1.1144e-13
C519 1612 2044 2.455e-14
C516 1615 2044 1.932e-14
C515 1616 2044 5.6e-14
C514 1617 2044 2.356e-14
C512 1619 2044 2.378e-14
C511 1620 2044 1.034e-13
C510 1621 2044 3.608e-14
C507 1624 2044 5.684e-14
C506 1625 2044 2.128e-14
C505 1626 2044 7.56e-15
C503 1628 2044 9.197e-14
C502 1629 2044 1.7149e-13
C500 1631 2044 1.853e-14
C499 1632 2044 9.81e-14
C498 1633 2044 6.05e-15
C497 1634 2044 5.123e-14
C496 1635 2044 1.8635e-14
C494 1637 2044 6.29e-14
C493 1638 2044 4.254e-14
C492 1639 2044 2.299e-14
C491 1640 2044 8.58e-15
C489 1642 2044 4.258e-14
C488 1643 2044 1.8635e-14
C487 1644 2044 6.05e-15
C486 1645 2044 4.867e-14
C484 1647 2044 1.853e-14
C483 1648 2044 4.922e-14
C481 1650 2044 2.299e-14
C480 1651 2044 1.2208e-13
C479 1652 2044 8.58e-15
C478 1653 2044 1.1718e-13
C477 1654 2044 4.3559e-13
C476 1655 2044 6.05e-15
C475 1656 2044 2.1957e-13
C474 1657 2044 9.5e-14
C473 1658 2044 1.8479e-13
C470 1661 2044 5.458e-14
C469 1662 2044 1.106e-13
C468 1663 2044 2.378e-14
C466 1665 2044 4.88e-14
C465 1666 2044 2.128e-14
C464 1667 2044 3.608e-14
C462 1669 2044 7.56e-15
C460 1671 2044 1.8635e-14
C458 1673 2044 6.3174e-13
C457 1674 2044 5.131e-14
C455 1676 2044 1.974e-13
C454 1677 2044 8.416e-14
C453 1678 2044 6.174e-14
C452 1679 2044 2.299e-14
C450 1681 2044 8.58e-15
C449 1682 2044 1.1815e-13
C448 1683 2044 4.686e-14
C447 1684 2044 9.678e-14
C446 1685 2044 5.218e-14
C445 1686 2044 1.8635e-14
C442 1689 2044 6.179e-14
C440 1691 2044 4.11e-15
C437 1694 2044 4.11e-15
C431 1700 2044 4.11e-15
C428 1703 2044 7.56e-15
C423 1708 2044 7.56e-15
C417 1714 2044 1.4934e-13
C416 1715 2044 6.05e-15
C414 1717 2044 6.05e-15
C412 1719 2044 6.05e-15
C410 1721 2044 8.68e-14
C408 1723 2044 8.58e-15
C406 1725 2044 4.11e-15
C399 1732 2044 6.05e-15
C396 1734 2044 9.7e-15
C395 1735 2044 1.0571e-13
C394 1736 2044 1.677e-14
C392 1738 2044 1.853e-14
C391 1739 2044 6.797e-14
C390 1740 2044 4.11e-15
C389 1741 2044 1.853e-14
C388 1742 2044 4.637e-14
C386 1744 2044 2.605e-14
C385 1745 2044 5.041e-14
C384 1746 2044 2.455e-14
C383 1747 2044 9.157e-14
C382 1748 2044 4.11e-15
C381 1749 2044 5.833e-14
C380 1750 2044 1.853e-14
C377 1753 2044 1.60938e-12
C376 1754 2044 5.477e-14
C375 1755 2044 7.883e-14
C373 1757 2044 5.4414e-13
C372 1758 2044 2.378e-14
C371 1759 2044 5.492e-14
C369 1761 2044 4.11e-15
C368 1762 2044 4.506e-14
C367 1763 2044 4.68e-14
C366 1764 2044 1.07117e-12
C365 1765 2044 2.212e-14
C362 1768 2044 7.56e-15
C361 1769 2044 1.3399e-13
C360 1770 2044 4.11e-15
C359 1771 2044 1.8635e-14
C358 1772 2044 6.4e-14
C357 1773 2044 2.378e-14
C355 1775 2044 2.128e-14
C354 1776 2044 5.208e-14
C353 1777 2044 7.56e-15
C350 1780 2044 3.608e-14
C347 1783 2044 5.507e-14
C346 1784 2044 5.578e-14
C345 1785 2044 4.11e-15
C344 1786 2044 2.455e-14
C342 1788 2044 1.767e-14
C341 1789 2044 1.6264e-13
C340 1790 2044 1.767e-14
C339 1791 2044 5.285e-14
C338 1792 2044 1.873e-13
C337 1793 2044 6.872e-14
C336 1794 2044 1.767e-14
C335 1795 2044 2.332e-13
C334 1796 2044 1.0488e-13
C333 1797 2044 2.299e-14
C332 1798 2044 4.11e-15
C331 1799 2044 1.8563e-13
C330 1800 2044 1.8635e-14
C328 1802 2044 4.258e-14
C327 1803 2044 1.8635e-14
C325 1805 2044 1.8635e-14
C323 1807 2044 7.268e-14
C322 1808 2044 1.8635e-14
C321 1809 2044 1.1148e-13
C319 1811 2044 4.11e-15
C318 1812 2044 5.233e-14
C316 1814 2044 2.605e-14
C315 1815 2044 4.11e-15
C314 1816 2044 1.0698e-13
C313 1817 2044 4.997e-14
C312 1818 2044 4.11e-15
C310 1820 2044 5.518e-14
C309 1821 2044 5.346e-14
C308 1822 2044 5.175e-14
C305 1825 2044 1.662e-14
C303 1827 2044 5.0667e-13
C300 1830 2044 1.8635e-14
C299 1831 2044 9.242e-14
C298 1832 2044 2.596e-14
C297 1833 2044 2.16e-14
C291 1838 2044 1.8635e-14
C290 1839 2044 6.453e-14
C288 1841 2044 1.853e-14
C287 1842 2044 1.316e-13
C286 1843 2044 4.763e-14
C285 1844 2044 6.05e-15
C282 1847 2044 2.455e-14
C281 1848 2044 8.237e-14
C280 1849 2044 1.19147e-12
C279 1850 2044 1.853e-14
C277 1852 2044 9.368e-14
C276 1853 2044 4.763e-14
C275 1854 2044 6.05e-15
C274 1855 2044 4.515e-14
C272 1857 2044 1.8635e-14
C271 1858 2044 9.077e-14
C269 1860 2044 5.057e-14
C266 1863 2044 1.853e-14
C265 1864 2044 1.9438e-13
C263 1866 2044 4.681e-14
C262 1867 2044 7.452e-14
C261 1868 2044 2.356e-14
C258 1871 2044 1.932e-14
C257 1872 2044 5e-14
C256 1873 2044 1.1946e-13
C255 1874 2044 1.8635e-14
C252 1877 2044 1.2806e-13
C251 1878 2044 1.095e-13
C250 1879 2044 1.8635e-14
C249 1880 2044 5.049e-14
C248 1881 2044 6.452e-14
C246 1883 2044 4.854e-14
C245 1884 2044 2.61056e-12
C244 1885 2044 8.678e-14
C243 1886 2044 4.877e-14
C242 1887 2044 1.767e-14
C241 1888 2044 6.05e-15
C240 1889 2044 1.767e-14
C239 1890 2044 6.05e-15
C238 1891 2044 1.1612e-13
C236 1893 2044 1.4111e-13
C235 1894 2044 1.8635e-14
C234 1895 2044 5.233e-14
C233 1896 2044 9.418e-14
C231 1898 2044 1.28652e-12
C230 1899 2044 1.41864e-12
C229 1900 2044 3.1404e-13
C228 1901 2044 8.805e-14
C227 1902 2044 5.061e-14
C226 1903 2044 6.547e-14
C224 1905 2044 6.05e-15
C223 1906 2044 1.8635e-14
C222 1907 2044 1.2206e-13
C221 1908 2044 2.596e-14
C220 1909 2044 2.16e-14
C219 1910 2044 7.76e-15
C213 1916 2044 9.7e-15
C208 1921 2044 6.05e-15
C207 1922 2044 7.76e-15
C205 1924 2044 7.76e-15
C202 1927 2044 7.76e-15
C201 1928 2044 6.05e-15
C198 1931 2044 6.05e-15
C195 1933 2044 2.659e-14
C194 1934 2044 1.568e-14
C193 1935 2044 1.0282e-13
C192 1936 2044 1.8635e-14
C190 1938 2044 1.677e-14
C189 1939 2044 4.11e-15
C188 1940 2044 4.963e-14
C187 1941 2044 7.277e-14
C186 1942 2044 1.853e-14
C184 1944 2044 4.11e-15
C182 1946 2044 1.8635e-14
C181 1947 2044 4.649e-14
C180 1948 2044 7.033e-14
C179 1949 2044 5.357e-14
C178 1950 2044 1.853e-14
C177 1951 2044 4.11e-15
C176 1952 2044 4.11e-15
C174 1954 2044 5.219e-14
C173 1955 2044 1.677e-14
C172 1956 2044 2.1408e-13
C170 1958 2044 1.8635e-14
C168 1960 2044 1.677e-14
C166 1962 2044 1.1298e-13
C165 1963 2044 2.596e-14
C162 1966 2044 1.2322e-13
C161 1967 2044 2.16e-14
C158 1970 2044 1.8635e-14
C156 1972 2044 7.757e-14
C155 1973 2044 5.281e-14
C154 1974 2044 1.853e-14
C153 1975 2044 4.11e-15
C152 1976 2044 5.057e-14
C151 1977 2044 2.9904e-13
C150 1978 2044 1.8635e-14
C149 1979 2044 7.43e-15
C148 1980 2044 1.662e-14
C147 1981 2044 2.3385e-13
C145 1983 2044 4.11e-15
C144 1984 2044 1.0819e-13
C143 1985 2044 1.677e-14
C140 1988 2044 1.0927e-13
C138 1990 2044 2.596e-14
C136 1992 2044 2.16e-14
C134 1994 2044 9.43e-14
C133 1995 2044 1.0102e-13
C131 1997 2044 1.8635e-14
C128 2000 2044 2.596e-14
C127 2001 2044 1.0454e-13
C126 2002 2044 2.16e-14
C122 2006 2044 1.8635e-14
C120 2008 2044 1.8635e-14
C118 2010 2044 1.2711e-13
C117 2011 2044 4.705e-14
C115 2013 2044 1.8635e-14
C114 2014 2044 1.2096e-13
C113 2015 2044 6.193e-14
C112 2016 2044 4.11e-15
C111 2017 2044 1.853e-14
C109 2019 2044 1.7631e-13
C108 2020 2044 2.596e-14
C106 2022 2044 1.4031e-13
C102 2026 2044 1.767e-14
C101 2027 2044 2.16e-14
C100 2028 2044 1.3082e-13
C99 2029 2044 9.236e-14
C98 2030 2044 4.541e-14
C95 2033 2044 1.8635e-14
C93 2035 2044 1.8635e-14
C92 2036 2044 1.1188e-13
C91 2037 2044 1.767e-14
C89 2039 2044 1.4096e-13
C87 2041 2044 8.446e-14
C86 2042 2044 1.8635e-14
C85 2043 2044 4.541e-14
C84 2044 2044 2.40799e-11
C83 2045 2044 7.253e-14
C82 2046 2044 1.677e-14
C80 2048 2044 4.963e-14
C79 2049 2044 4.649e-14
C78 2050 2044 1.853e-14
C76 2052 2044 1.677e-14
C74 2054 2044 1.8635e-14
C73 2055 2044 2.6736e-12
C72 2056 2044 1.0469e-13
C71 2057 2044 1.853e-14
C70 2058 2044 4.22515e-12
C69 2059 2044 4.963e-14
C68 2060 2044 1.8635e-14
C66 2062 2044 4.649e-14
C65 2063 2044 1.0866e-13
C64 2064 2044 1.8635e-14
C63 2065 2044 2.596e-14
C62 2066 2044 1.0104e-13
C61 2067 2044 2.16e-14
C60 2068 2044 7.76e-15
C59 2069 2044 1.1242e-13
C58 2070 2044 1.4466e-13
C57 2071 2044 1.8635e-14
C56 2072 2044 1.8635e-14
C54 2074 2044 2.1747e-13
C53 2075 2044 8.666e-14
C50 2078 2044 2.639e-14
C49 2079 2044 1.0758e-13
C48 2080 2044 1.853e-14
C46 2082 2044 2.596e-14
C45 2083 2044 8.576e-14
C44 2084 2044 2.16e-14
C43 2085 2044 7.76e-15
C41 2087 2044 8.982e-14
C40 2088 2044 4.361e-13
C39 2089 2044 1.568e-14
C38 2090 2044 1.8635e-14
C36 2092 2044 1.4499e-13
C35 2093 2044 2.1231e-13
C34 2094 2044 6.05e-15
C33 2095 2044 5.157e-14
C32 2096 2044 3.1681e-13
C31 2097 2044 2.596e-14
C30 2098 2044 1.3706e-13
C29 2099 2044 9.7e-15
C28 2100 2044 2.16e-14
C27 2101 2044 2.3098e-13
C26 2102 2044 8.912e-14
C25 2103 2044 1.568e-14
C24 2104 2044 1.4223e-13
C23 2105 2044 1.96016e-12
C21 2107 2044 1.8635e-14
C20 2108 2044 3.24469e-12
C19 2109 2044 1.6647e-13
C18 2110 2044 2.596e-14
C17 2111 2044 2.1461e-13
C16 2112 2044 7.76e-15
C15 2113 2044 3.53277e-12
C14 2114 2044 2.16e-14
C13 2115 2044 1.71672e-12
C12 2116 2044 2.596e-14
C11 2117 2044 2.16e-14
C10 2118 2044 7.76e-15
C9 2119 2044 8.878e-14
C8 2120 2044 8.34e-14
C7 2121 2044 1.0546e-13
C6 2122 2044 1.73654e-12
C5 2123 2044 1.4815e-12
C4 2124 2044 1.8635e-14
C3 2125 2044 1.96098e-12
C2 2126 2044 1.45569e-12
C1 2127 2044 2.49659e-11
.ends mul5b_cougar

