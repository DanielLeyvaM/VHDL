* Spice description of sum2b_cougar
* Spice driver version -1209303388
* Date ( dd/mm/yyyy hh:mm:ss ): 28/10/2020 at 12:54:11

* INTERF a[0] a[1] b[0] b[1] ci co so[0] so[1] vdd vss 


.subckt sum2b_cougar 24 39 8 40 9 37 26 17 44 30 
* NET 8 = b[0]
* NET 9 = ci
* NET 17 = so[1]
* NET 24 = a[0]
* NET 25 = xr2_x1_sig
* NET 26 = so[0]
* NET 30 = vss
* NET 33 = xr2_x1_2_sig
* NET 37 = co
* NET 38 = aux3
* NET 39 = a[1]
* NET 40 = b[1]
* NET 41 = a2_x2_sig
* NET 44 = vdd
Mtr_00076 41 36 44 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00075 44 39 36 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 36 40 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 45 38 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 43 39 42 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 44 40 43 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 42 41 45 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 37 42 44 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00068 32 40 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 44 39 35 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 33 32 34 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00065 34 39 44 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00064 34 35 33 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00063 44 40 34 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00062 23 24 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 44 25 28 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 26 23 14 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00059 14 25 44 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00058 14 28 26 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00057 44 24 14 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00056 15 33 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 44 38 19 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 17 15 13 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00053 13 38 44 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00052 13 19 17 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00051 44 33 13 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00050 10 8 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 44 9 12 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 25 10 11 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00047 11 9 44 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00046 11 12 25 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00045 44 8 11 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00044 38 5 44 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00043 7 9 6 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00042 7 8 44 44 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00041 44 9 7 44 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00040 6 8 5 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00039 5 24 7 44 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00038 36 40 22 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 30 36 41 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 22 39 30 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 31 39 30 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 30 40 31 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 31 38 42 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 42 41 31 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00031 30 42 37 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 35 39 30 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 30 40 32 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 16 32 30 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 33 35 16 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 21 40 33 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 30 39 21 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 28 25 30 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 30 24 23 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 29 23 30 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 26 28 29 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 27 24 26 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 30 25 27 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 19 38 30 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 30 33 15 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 20 15 30 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 17 19 20 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 18 33 17 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 30 38 18 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 12 9 30 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 30 8 10 30 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 4 10 30 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 25 12 4 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 3 8 25 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 30 9 3 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 30 5 38 30 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 30 8 2 30 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00004 2 9 30 30 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00003 5 8 1 30 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00002 1 9 30 30 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00001 2 24 5 30 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
C46 2 30 4.11e-15
C42 5 30 2.299e-14
C40 7 30 8.58e-15
C39 8 30 9.68e-14
C38 9 30 9.907e-14
C37 10 30 2.596e-14
C36 11 30 9.7e-15
C35 12 30 2.16e-14
C34 13 30 9.7e-15
C32 14 30 9.7e-15
C31 15 30 2.596e-14
C29 17 30 3.889e-14
C27 19 30 2.16e-14
C23 23 30 2.596e-14
C22 24 30 8.045e-14
C21 25 30 5.991e-14
C20 26 30 5.905e-14
C18 28 30 2.16e-14
C16 30 30 4.2076e-13
C15 31 30 7.43e-15
C14 32 30 2.596e-14
C13 33 30 6.235e-14
C12 34 30 9.7e-15
C11 35 30 2.16e-14
C10 36 30 1.8635e-14
C9 37 30 3.288e-14
C8 38 30 1.185e-13
C7 39 30 1.0297e-13
C6 40 30 1.0289e-13
C5 41 30 5.503e-14
C4 42 30 2.639e-14
C2 44 30 4.2692e-13
.ends sum2b_cougar

