* Spice description of sum4b_cougar
* Spice driver version -1208795484
* Date ( dd/mm/yyyy hh:mm:ss ): 26/10/2020 at 21:04:52

* INTERF a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] ci co so[0] so[1] so[2] 
* INTERF so[3] vdd vss 


.subckt sum4b_cougar 132 121 88 52 130 119 113 114 131 7 116 108 76 34 136 106 
* NET 5 = inv_x2_2_sig
* NET 7 = co
* NET 9 = o3_x2_sig
* NET 12 = o4_x2_sig
* NET 16 = inv_x2_sig
* NET 17 = o2_x2_sig
* NET 20 = aux0
* NET 26 = inv_x2_3_sig
* NET 27 = mbk_buf_aux12
* NET 30 = na3_x1_sig
* NET 34 = so[3]
* NET 35 = not_aux13
* NET 36 = aux7
* NET 39 = na4_x1_sig
* NET 41 = na4_x1_2_sig
* NET 42 = na2_x1_2_sig
* NET 52 = a[3]
* NET 56 = aux12
* NET 58 = not_aux11
* NET 60 = mbk_buf_not_aux11
* NET 61 = aux13
* NET 62 = not_b[2]
* NET 63 = na2_x1_sig
* NET 64 = not_aux5
* NET 65 = na3_x1_2_sig
* NET 67 = aux5
* NET 68 = not_a[1]
* NET 76 = so[2]
* NET 81 = mbk_buf_aux11
* NET 82 = xr2_x1_3_sig
* NET 88 = a[2]
* NET 90 = aux11
* NET 95 = a2_x2_sig
* NET 100 = aux6
* NET 102 = not_b[1]
* NET 103 = not_aux4
* NET 106 = vss
* NET 108 = so[1]
* NET 112 = mbk_buf_aux4
* NET 113 = b[2]
* NET 114 = b[3]
* NET 116 = so[0]
* NET 119 = b[1]
* NET 121 = a[1]
* NET 123 = xr2_x1_2_sig
* NET 126 = xr2_x1_sig
* NET 128 = aux4
* NET 130 = b[0]
* NET 131 = ci
* NET 132 = a[0]
* NET 136 = vdd
Mtr_00252 128 133 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00251 135 130 134 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00250 135 131 136 136 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00249 136 130 135 136 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00248 134 131 133 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00247 133 132 135 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00246 125 131 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00245 136 130 129 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 126 125 127 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00243 127 130 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00242 127 129 126 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00241 136 131 127 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00240 112 110 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00239 136 128 110 136 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00238 120 119 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 136 121 124 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 123 120 122 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00235 122 121 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00234 122 124 123 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00233 136 119 122 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00232 107 123 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 136 112 111 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 108 107 109 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00229 109 112 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00228 109 111 108 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00227 136 123 109 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00226 115 132 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00225 136 126 118 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00224 116 115 117 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00223 117 126 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00222 117 118 116 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00221 136 132 117 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00220 95 97 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00219 136 121 97 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 97 119 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 100 102 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 136 103 100 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00215 103 128 136 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00214 72 128 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 71 121 92 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 136 119 71 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 92 95 72 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00210 90 92 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00209 102 119 136 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00208 84 113 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 136 88 89 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 82 84 70 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00205 70 88 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00204 70 89 82 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00203 136 113 70 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00202 73 82 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 136 81 80 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 76 73 69 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00199 69 81 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00198 69 80 76 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00197 136 82 69 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00196 81 79 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00195 136 90 79 136 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00194 66 103 67 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00193 136 102 66 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00192 64 67 136 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00191 68 121 136 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00190 63 62 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00189 136 60 63 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00188 136 63 65 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00187 65 61 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00186 65 88 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00185 62 113 136 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00184 136 90 58 136 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_00183 58 90 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00182 60 59 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00181 136 58 59 136 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00180 55 58 57 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00179 136 62 55 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00178 56 57 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00177 136 50 24 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00176 24 51 61 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00175 24 52 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00174 61 114 24 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00173 136 52 51 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00172 50 114 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 136 100 36 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 36 47 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 136 68 47 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 42 68 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 136 64 42 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 136 113 41 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00165 41 42 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00164 136 61 41 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00163 41 100 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 136 62 39 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 39 35 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00160 136 36 39 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 39 64 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 35 61 136 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00157 136 35 30 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00156 30 27 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00155 30 26 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 27 25 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00153 136 56 25 136 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00152 136 41 34 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 34 39 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 136 30 34 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 34 65 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00148 20 21 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00147 136 114 21 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 21 52 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00145 16 36 136 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00144 19 114 18 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00143 136 52 19 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00142 17 18 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00141 14 16 13 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00140 15 113 14 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00139 11 20 15 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00138 136 67 11 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00137 136 13 12 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00136 136 88 4 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00135 4 20 8 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00134 8 5 6 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00133 9 6 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00132 136 9 10 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00131 7 10 136 136 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00130 136 17 10 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 10 12 136 136 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 26 88 136 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00127 5 56 136 136 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00126 106 133 128 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 106 131 105 106 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00124 105 130 106 106 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00123 133 131 104 106 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00122 104 130 106 106 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00121 105 132 133 106 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00120 129 130 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00119 106 131 125 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00118 98 125 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 126 129 98 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 99 131 126 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 106 130 99 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 106 110 112 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 110 128 106 106 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00112 124 121 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00111 106 119 120 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00110 91 120 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 123 124 91 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 93 119 123 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00107 106 121 93 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 111 112 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00105 106 123 107 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00104 78 107 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 108 111 78 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 77 123 108 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 106 112 77 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 118 126 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00099 106 132 115 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00098 87 115 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 116 118 87 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 86 132 116 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 106 126 86 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 97 119 96 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 106 97 95 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00092 96 121 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 106 102 101 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 101 103 100 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 106 128 103 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 94 121 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00087 106 119 94 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00086 94 128 92 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00085 92 95 94 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00084 106 92 90 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 106 119 102 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 89 88 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00081 106 113 84 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00080 85 84 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 82 89 85 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 83 113 82 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 106 88 83 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 80 81 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00075 106 82 73 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00074 75 73 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 76 80 75 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 74 82 76 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 106 81 74 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 106 79 81 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 79 90 106 106 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00068 67 102 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00067 106 103 67 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00066 106 67 64 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 106 121 68 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 106 62 46 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 46 60 63 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 106 88 49 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 49 63 48 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 48 61 65 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 106 113 62 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 106 90 58 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 58 90 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 106 59 60 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 59 58 106 106 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00054 56 57 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 57 62 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00052 106 58 57 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00051 106 52 54 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 54 50 61 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 61 51 53 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 53 114 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 106 114 50 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 51 52 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 47 68 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00044 23 100 36 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 106 47 23 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 106 68 22 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 22 64 42 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 106 100 45 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 45 113 44 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 44 42 43 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 43 61 41 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 106 64 40 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 40 62 37 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 37 35 38 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 38 36 39 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 106 61 35 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 106 26 29 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 29 35 28 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 28 27 30 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 106 25 27 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 25 56 106 106 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00026 106 65 31 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 31 41 33 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 33 39 32 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 32 30 34 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 21 52 3 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 106 21 20 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 3 114 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 106 36 16 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 17 18 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 18 52 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 106 114 18 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 13 67 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 106 16 13 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 106 20 13 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 13 113 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 12 13 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 6 5 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 6 88 106 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 106 20 6 106 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 106 6 9 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 106 10 7 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 2 9 106 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 1 12 2 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 10 17 1 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 106 88 26 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 106 56 5 106 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C135 5 106 5.619e-14
C134 6 106 2.455e-14
C133 7 106 4.016e-14
C131 9 106 5.627e-14
C130 10 106 2.605e-14
C128 12 106 4.909e-14
C127 13 106 2.72e-14
C124 16 106 4.419e-14
C123 17 106 6.071e-14
C122 18 106 1.8635e-14
C120 20 106 1.0064e-13
C119 21 106 1.8635e-14
C115 24 106 7.76e-15
C114 25 106 1.568e-14
C113 26 106 5.759e-14
C112 27 106 5.008e-14
C109 30 106 5.64e-14
C105 34 106 4.715e-14
C104 35 106 8.84e-14
C103 36 106 1.0437e-13
C100 39 106 5.396e-14
C98 41 106 6.266e-14
C97 42 106 5.166e-14
C92 47 106 1.662e-14
C89 50 106 2.596e-14
C88 51 106 2.16e-14
C87 52 106 9.176e-14
C82 56 106 9.004e-14
C81 57 106 1.8635e-14
C80 58 106 7.858e-14
C79 59 106 1.568e-14
C78 60 106 5.838e-14
C77 61 106 1.3603e-13
C76 62 106 1.3612e-13
C75 63 106 5.566e-14
C74 64 106 1.0614e-13
C73 65 106 7.92e-14
C71 67 106 1.0942e-13
C70 68 106 1.0022e-13
C69 69 106 9.7e-15
C68 70 106 9.7e-15
C64 73 106 2.596e-14
C61 76 106 5.185e-14
C58 79 106 1.568e-14
C57 80 106 2.16e-14
C56 81 106 5.169e-14
C55 82 106 7.435e-14
C53 84 106 2.596e-14
C49 88 106 2.1523e-13
C48 89 106 2.16e-14
C47 90 106 1.0138e-13
C45 92 106 2.639e-14
C43 94 106 7.43e-15
C42 95 106 4.783e-14
C40 97 106 1.8635e-14
C37 100 106 1.152e-13
C35 102 106 8.715e-14
C34 103 106 8.1e-14
C32 105 106 4.11e-15
C31 106 106 1.47812e-12
C30 107 106 2.596e-14
C29 108 106 4.249e-14
C28 109 106 9.7e-15
C27 110 106 1.568e-14
C26 111 106 2.16e-14
C25 112 106 5.169e-14
C24 113 106 1.8231e-13
C23 114 106 1.8939e-13
C22 115 106 2.596e-14
C21 116 106 4.681e-14
C20 117 106 9.7e-15
C19 118 106 2.16e-14
C18 119 106 1.3724e-13
C17 120 106 2.596e-14
C16 121 106 1.5687e-13
C15 122 106 9.7e-15
C14 123 106 8.395e-14
C13 124 106 2.16e-14
C12 125 106 2.596e-14
C11 126 106 6.831e-14
C10 127 106 9.7e-15
C9 128 106 1.6881e-13
C8 129 106 2.16e-14
C7 130 106 8.675e-14
C6 131 106 1.416e-13
C5 132 106 9.6e-14
C4 133 106 2.299e-14
C2 135 106 8.58e-15
C1 136 106 1.54056e-12
.ends sum4b_cougar

