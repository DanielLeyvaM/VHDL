* Spice description of sum3b_cougar
* Spice driver version -1208856924
* Date ( dd/mm/yyyy hh:mm:ss ):  9/10/2020 at 20:39:58

* INTERF a[0] a[1] a[2] b[0] b[1] b[2] ci co so[0] so[1] so[2] vdd vss 


.subckt sum3b_cougar a[0] a[1] a[2] b[0] b[1] b[2] ci co so[0] so[1] so[2] vdd vss 
Mtr_00118 acarreo0 sig4 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00117 sig2 cix sig3 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00116 sig2 a[0] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00115 vdd cix sig2 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00114 sig3 a[0] sig4 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00113 sig4 b[0] sig2 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00112 sig12 a[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 vdd cix sig9 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 x0.xr2_x1_sig sig12 sig10 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00109 sig10 cix vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00108 sig10 sig9 x0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00107 vdd a[0] sig10 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00106 sig17 b[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 vdd x0.xr2_x1_sig sig16 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 so[0] sig17 sig14 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00103 sig14 x0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00102 sig14 sig16 so[0] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00101 vdd b[0] sig14 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00100 acarreo1 sig28 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00099 sig49 acarreo0 sig50 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00098 sig49 a[1] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00097 vdd acarreo0 sig49 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00096 sig50 a[1] sig28 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00095 sig28 b[1] sig49 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00094 sig26 a[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 vdd acarreo0 sig23 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00092 x1.xr2_x1_sig sig26 sig47 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00091 sig47 acarreo0 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00090 sig47 sig23 x1.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00089 vdd a[1] sig47 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00088 sig45 b[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 vdd x2.xr2_x1_sig sig42 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 so[2] sig45 sig52 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00085 sig52 x2.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00084 sig52 sig42 so[2] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00083 vdd b[2] sig52 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00082 sig38 b[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 vdd x1.xr2_x1_sig sig33 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 so[1] sig38 sig51 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00079 sig51 x1.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00078 sig51 sig33 so[1] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00077 vdd b[1] sig51 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00076 vdd ci sig53 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00075 vdd sig53 cix vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00074 cix sig53 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00073 vdd sig53 cix vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00072 cix sig53 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00071 sig58 a[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 vdd acarreo1 sig56 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 x2.xr2_x1_sig sig58 sig57 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00068 sig57 acarreo1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00067 sig57 sig56 x2.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00066 vdd a[2] sig57 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00065 co sig61 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00064 sig59 acarreo1 sig60 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00063 sig59 a[2] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00062 vdd acarreo1 sig59 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00061 sig60 a[2] sig61 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00060 sig61 b[2] sig59 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00059 vss sig4 acarreo0 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 vss a[0] sig19 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00057 sig19 cix vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00056 sig4 a[0] sig21 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00055 sig21 cix vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00054 sig19 b[0] sig4 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00053 sig9 cix vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00052 vss a[0] sig12 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00051 sig34 sig12 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 x0.xr2_x1_sig sig9 sig34 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 sig30 a[0] x0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 vss cix sig30 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 sig16 x0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 vss b[0] sig17 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 sig40 sig17 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 so[0] sig16 sig40 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 sig39 b[0] so[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 vss x0.xr2_x1_sig sig39 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 vss sig28 acarreo1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 vss a[1] sig32 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00039 sig32 acarreo0 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00038 sig28 a[1] sig29 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00037 sig29 acarreo0 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00036 sig32 b[1] sig28 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00035 sig23 acarreo0 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 vss a[1] sig26 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 sig22 sig26 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 x1.xr2_x1_sig sig23 sig22 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 sig24 a[1] x1.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 vss acarreo0 sig24 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 sig42 x2.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 vss b[2] sig45 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00027 sig46 sig45 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 so[2] sig42 sig46 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 sig41 b[2] so[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 vss x2.xr2_x1_sig sig41 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 sig33 x1.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 vss b[1] sig38 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00021 sig37 sig38 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 so[1] sig33 sig37 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 sig35 b[1] so[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 vss x1.xr2_x1_sig sig35 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 sig53 ci vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 cix sig53 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 vss sig53 cix vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 vss sig53 cix vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 cix sig53 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 sig56 acarreo1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 vss a[2] sig58 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 sig65 sig58 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 x2.xr2_x1_sig sig56 sig65 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 sig64 a[2] x2.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 vss acarreo1 sig64 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 vss sig61 co vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 vss a[2] sig66 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00004 sig66 acarreo1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00003 sig61 a[2] sig67 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00002 sig67 acarreo1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00001 sig66 b[2] sig61 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
C66 sig66 vss 4.11e-15
C62 co vss 3.8e-14
C61 sig61 vss 2.299e-14
C59 sig59 vss 8.58e-15
C58 sig58 vss 2.596e-14
C57 sig57 vss 9.7e-15
C56 sig56 vss 2.16e-14
C55 a[2] vss 1.0123e-13
C54 ci vss 4.245e-14
C53 sig53 vss 4.103e-14
C52 sig52 vss 9.7e-15
C51 sig51 vss 9.7e-15
C49 sig49 vss 8.58e-15
C47 sig47 vss 9.7e-15
C45 sig45 vss 2.596e-14
C44 so[2] vss 4.009e-14
C43 x2.xr2_x1_sig vss 7.431e-14
C42 sig42 vss 2.16e-14
C38 sig38 vss 2.596e-14
C36 so[1] vss 4.489e-14
C33 sig33 vss 2.16e-14
C32 sig32 vss 4.11e-15
C31 acarreo1 vss 1.2771e-13
C28 sig28 vss 2.299e-14
C27 a[1] vss 8.491e-14
C26 sig26 vss 2.596e-14
C25 x1.xr2_x1_sig vss 6.951e-14
C23 sig23 vss 2.16e-14
C20 vss vss 6.43161e-13
C19 sig19 vss 4.11e-15
C18 b[2] vss 9.485e-14
C17 sig17 vss 2.596e-14
C16 sig16 vss 2.16e-14
C15 so[0] vss 3.649e-14
C14 sig14 vss 9.7e-15
C13 b[1] vss 8.621e-14
C12 sig12 vss 2.596e-14
C11 x0.xr2_x1_sig vss 6.111e-14
C10 sig10 vss 9.7e-15
C9 sig9 vss 2.16e-14
C8 acarreo0 vss 1.0627e-13
C7 cix vss 1.3659e-13
C6 a[0] vss 9.211e-14
C5 b[0] vss 9.725e-14
C4 sig4 vss 2.299e-14
C2 sig2 vss 8.58e-15
C1 vdd vss 6.52121e-13
.ends sum3b_cougar

