* Spice description of mux41_cougar
* Spice driver version -1208709468
* Date ( dd/mm/yyyy hh:mm:ss ): 28/09/2020 at 18:40:59

* INTERF a b c d s[0] s[1] vdd vss x 


.subckt mux41_cougar 11 5 25 16 20 26 30 13 15 
* NET 5 = b
* NET 7 = on12_x1_2_sig
* NET 11 = a
* NET 12 = not_s[1]
* NET 13 = vss
* NET 14 = na3_x1_sig
* NET 15 = x
* NET 16 = d
* NET 18 = on12_x1_sig
* NET 19 = an12_x1_sig
* NET 20 = s[0]
* NET 21 = o3_x2_sig
* NET 25 = c
* NET 26 = s[1]
* NET 28 = an12_x1_2_sig
* NET 30 = vdd
Mtr_00050 30 20 24 30 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00049 24 28 22 30 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00048 22 19 23 30 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00047 21 23 30 30 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00046 27 26 30 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 30 27 29 30 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00044 29 25 28 30 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00043 15 14 30 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 30 21 15 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 30 26 18 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 18 17 30 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 30 16 17 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 12 26 30 30 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00037 30 26 12 30 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00036 30 26 12 30 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00035 12 26 30 30 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00034 10 12 30 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 30 10 1 30 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00032 1 11 19 30 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00031 30 12 7 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 7 6 30 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 30 5 6 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 30 20 14 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 14 18 30 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 14 7 30 30 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 23 19 13 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00024 23 20 13 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 13 28 23 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 13 23 21 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 13 26 27 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 28 27 13 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00019 13 25 28 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 13 14 4 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 4 21 15 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 17 16 13 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 9 26 18 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 13 17 9 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 13 26 12 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 12 26 13 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 13 26 12 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 12 26 13 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 13 12 10 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 19 10 13 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 13 11 19 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 6 5 13 13 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 8 12 7 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 13 6 8 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 13 7 2 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 2 20 3 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 3 18 14 13 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C26 5 13 3.429e-14
C25 6 13 1.662e-14
C24 7 13 5.201e-14
C21 10 13 1.677e-14
C20 11 13 3.736e-14
C19 12 13 1.0759e-13
C18 13 13 2.8924e-13
C17 14 13 6.113e-14
C16 15 13 2.757e-14
C15 16 13 3.429e-14
C14 17 13 1.662e-14
C13 18 13 5.994e-14
C12 19 13 5.221e-14
C11 20 13 7.732e-14
C10 21 13 6.202e-14
C8 23 13 2.455e-14
C6 25 13 3.52e-14
C5 26 13 1.5361e-13
C4 27 13 1.677e-14
C3 28 13 5.143e-14
C1 30 13 2.9904e-13
.ends mux41_cougar

