* Spice description of sum5b_cougar
* Spice driver version -1209602396
* Date ( dd/mm/yyyy hh:mm:ss ): 28/10/2020 at 12:59:36

* INTERF a[0] a[1] a[2] a[3] a[4] b[0] b[1] b[2] b[3] b[4] ci co so[0] so[1] 
* INTERF so[2] so[3] so[4] vdd vss 


.subckt sum5b_cougar a[0] a[1] a[2] a[3] a[4] b[0] b[1] b[2] b[3] b[4] ci co so[0] so[1] so[2] so[3] so[4] vdd vss 
Mtr_00190 acarreo0 sig4 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00189 sig2 cix sig3 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00188 sig2 b[0] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00187 vdd cix sig2 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00186 sig3 b[0] sig4 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00185 sig4 a[0] sig2 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00184 sig18 b[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 vdd cix sig14 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00182 x0.xr2_x1_sig sig18 sig15 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00181 sig15 cix vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00180 sig15 sig14 x0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00179 vdd b[0] sig15 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00178 sig23 a[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00177 vdd x0.xr2_x1_sig sig20 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 so[0] sig23 sig21 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00175 sig21 x0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00174 sig21 sig20 so[0] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00173 vdd a[0] sig21 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00172 sig12 b[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 vdd acarreo0 sig8 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 x1.xr2_x1_sig sig12 sig10 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00169 sig10 acarreo0 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00168 sig10 sig8 x1.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00167 vdd b[1] sig10 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00166 acarreo2 sig36 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00165 sig57 acarreo1 sig58 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00164 sig57 b[2] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00163 vdd acarreo1 sig57 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00162 sig58 b[2] sig36 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00161 sig36 a[2] sig57 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00160 acarreo1 sig29 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00159 sig55 acarreo0 sig56 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00158 sig55 b[1] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00157 vdd acarreo0 sig55 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00156 sig56 b[1] sig29 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00155 sig29 a[1] sig55 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00154 sig53 b[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00153 vdd acarreo2 sig49 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 x3.xr2_x1_sig sig53 sig60 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00151 sig60 acarreo2 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00150 sig60 sig49 x3.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00149 vdd b[3] sig60 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00148 sig44 a[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 vdd x1.xr2_x1_sig sig40 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 so[1] sig44 sig59 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00145 sig59 x1.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00144 sig59 sig40 so[1] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00143 vdd a[1] sig59 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00142 sig68 b[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 vdd acarreo1 sig67 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 x2.xr2_x1_sig sig68 sig69 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00139 sig69 acarreo1 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00138 sig69 sig67 x2.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00137 vdd b[2] sig69 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00136 sig64 a[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 vdd x2.xr2_x1_sig sig61 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 so[2] sig64 sig62 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00133 sig62 x2.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00132 sig62 sig61 so[2] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00131 vdd a[2] sig62 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00130 sig77 a[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 vdd x3.xr2_x1_sig sig74 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 so[3] sig77 sig76 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00127 sig76 x3.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00126 sig76 sig74 so[3] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00125 vdd a[3] sig76 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00124 acarreo3 sig73 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00123 sig70 acarreo2 sig71 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00122 sig70 b[3] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00121 vdd acarreo2 sig70 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00120 sig71 b[3] sig73 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00119 sig73 a[3] sig70 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00118 sig91 a[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 vdd x4.xr2_x1_sig sig90 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 so[4] sig91 sig102 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00115 sig102 x4.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00114 sig102 sig90 so[4] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00113 vdd a[4] sig102 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00112 vdd ci sig81 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00111 vdd sig81 cix vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00110 cix sig81 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00109 vdd sig81 cix vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00108 cix sig81 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00107 sig97 b[4] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 vdd acarreo3 sig96 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 x4.xr2_x1_sig sig97 sig103 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00104 sig103 acarreo3 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00103 sig103 sig96 x4.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00102 vdd b[4] sig103 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00101 co sig100 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00100 sig106 acarreo3 sig107 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00099 sig106 b[4] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00098 vdd acarreo3 sig106 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00097 sig107 b[4] sig100 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00096 sig100 a[4] sig106 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00095 vss sig4 acarreo0 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 vss b[0] sig26 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00093 sig26 cix vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00092 sig4 b[0] sig28 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00091 sig28 cix vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00090 sig26 a[0] sig4 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00089 sig14 cix vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00088 vss b[0] sig18 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00087 sig42 sig18 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 x0.xr2_x1_sig sig14 sig42 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 sig39 b[0] x0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00084 vss cix sig39 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 sig20 x0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00082 vss a[0] sig23 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00081 sig51 sig23 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 so[0] sig20 sig51 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 sig47 a[0] so[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 vss x0.xr2_x1_sig sig47 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 sig8 acarreo0 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00076 vss b[1] sig12 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00075 sig33 sig12 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 x1.xr2_x1_sig sig8 sig33 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 sig34 b[1] x1.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 vss acarreo0 sig34 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 vss sig36 acarreo2 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 vss b[2] sig35 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00069 sig35 acarreo1 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00068 sig36 b[2] sig37 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00067 sig37 acarreo1 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00066 sig35 a[2] sig36 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00065 vss sig29 acarreo1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 vss b[1] sig27 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00063 sig27 acarreo0 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00062 sig29 b[1] sig30 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00061 sig30 acarreo0 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00060 sig27 a[1] sig29 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00059 sig49 acarreo2 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00058 vss b[3] sig53 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00057 sig52 sig53 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 x3.xr2_x1_sig sig49 sig52 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 sig50 b[3] x3.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 vss acarreo2 sig50 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 sig40 x1.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00052 vss a[1] sig44 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00051 sig43 sig44 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 so[1] sig40 sig43 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 sig45 a[1] so[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 vss x1.xr2_x1_sig sig45 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 sig67 acarreo1 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 vss b[2] sig68 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 sig84 sig68 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 x2.xr2_x1_sig sig67 sig84 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 sig85 b[2] x2.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 vss acarreo1 sig85 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 sig61 x2.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00040 vss a[2] sig64 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00039 sig80 sig64 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 so[2] sig61 sig80 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 sig79 a[2] so[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 vss x2.xr2_x1_sig sig79 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 sig74 x3.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 vss a[3] sig77 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 sig99 sig77 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 so[3] sig74 sig99 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 sig98 a[3] so[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 vss x3.xr2_x1_sig sig98 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 vss sig73 acarreo3 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 vss b[3] sig94 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00027 sig94 acarreo2 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00026 sig73 b[3] sig93 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00025 sig93 acarreo2 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00024 sig94 a[3] sig73 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00023 sig90 x4.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 vss a[4] sig91 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00021 sig88 sig91 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 so[4] sig90 sig88 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 sig86 a[4] so[4] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 vss x4.xr2_x1_sig sig86 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 sig81 ci vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 cix sig81 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 vss sig81 cix vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 vss sig81 cix vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 cix sig81 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 sig96 acarreo3 vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 vss b[4] sig97 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 sig95 sig97 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 x4.xr2_x1_sig sig96 sig95 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 sig92 b[4] x4.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 vss acarreo3 sig92 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 vss sig100 co vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 vss b[4] sig104 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00004 sig104 acarreo3 vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00003 sig100 b[4] sig105 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00002 sig105 acarreo3 vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00001 sig104 a[4] sig100 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
C108 co vss 3.92e-14
C106 sig106 vss 8.58e-15
C104 sig104 vss 4.11e-15
C103 sig103 vss 9.7e-15
C102 sig102 vss 9.7e-15
C100 sig100 vss 2.299e-14
C97 sig97 vss 2.596e-14
C96 sig96 vss 2.16e-14
C94 sig94 vss 4.11e-15
C91 sig91 vss 2.596e-14
C90 sig90 vss 2.16e-14
C89 a[4] vss 9.36e-14
C87 so[4] vss 6.001e-14
C83 x4.xr2_x1_sig vss 6.351e-14
C82 ci vss 4.485e-14
C81 sig81 vss 4.103e-14
C77 sig77 vss 2.596e-14
C76 sig76 vss 9.7e-15
C75 so[3] vss 3.241e-14
C74 sig74 vss 2.16e-14
C73 sig73 vss 2.299e-14
C72 acarreo3 vss 1.1155e-13
C70 sig70 vss 8.58e-15
C69 sig69 vss 9.7e-15
C68 sig68 vss 2.596e-14
C67 sig67 vss 2.16e-14
C66 a[3] vss 1.044e-13
C65 x2.xr2_x1_sig vss 6.351e-14
C64 sig64 vss 2.596e-14
C63 so[2] vss 8.089e-14
C62 sig62 vss 9.7e-15
C61 sig61 vss 2.16e-14
C60 sig60 vss 9.7e-15
C59 sig59 vss 9.7e-15
C57 sig57 vss 8.58e-15
C55 sig55 vss 8.58e-15
C53 sig53 vss 2.596e-14
C49 sig49 vss 2.16e-14
C48 x3.xr2_x1_sig vss 5.991e-14
C46 so[1] vss 4.321e-14
C44 sig44 vss 2.596e-14
C41 acarreo2 vss 1.1755e-13
C40 sig40 vss 2.16e-14
C38 a[2] vss 8.208e-14
C36 sig36 vss 2.299e-14
C35 sig35 vss 4.11e-15
C32 acarreo1 vss 1.0563e-13
C31 a[1] vss 9.888e-14
C29 sig29 vss 2.299e-14
C27 sig27 vss 4.11e-15
C26 sig26 vss 4.11e-15
C25 vss vss 1.00728e-12
C24 b[4] vss 1.212e-13
C23 sig23 vss 2.596e-14
C22 so[0] vss 3.241e-14
C21 sig21 vss 9.7e-15
C20 sig20 vss 2.16e-14
C19 b[3] vss 1.2672e-13
C18 sig18 vss 2.596e-14
C17 b[2] vss 1.1576e-13
C16 x0.xr2_x1_sig vss 5.991e-14
C15 sig15 vss 9.7e-15
C14 sig14 vss 2.16e-14
C13 b[1] vss 1.0968e-13
C12 sig12 vss 2.596e-14
C11 x1.xr2_x1_sig vss 6.831e-14
C10 sig10 vss 9.7e-15
C9 acarreo0 vss 1.1275e-13
C8 sig8 vss 2.16e-14
C7 cix vss 1.5819e-13
C6 b[0] vss 1.0392e-13
C5 a[0] vss 9.96e-14
C4 sig4 vss 2.299e-14
C2 sig2 vss 8.58e-15
C1 vdd vss 1.01456e-12
.ends sum5b_cougar

