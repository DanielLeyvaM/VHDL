* Spice description of mul3b_cougar
* Spice driver version -1209459036
* Date ( dd/mm/yyyy hh:mm:ss ): 28/10/2020 at 14:33:46

* INTERF vdd vss x[0] x[1] x[2] y[0] y[1] y[2] z[0] z[1] z[2] z[3] z[4] z[5] 


.subckt mul3b_cougar 167 140 156 158 163 149 164 131 141 143 74 54 27 3 
* NET 3 = z[5]
* NET 6 = an12_x1_sig
* NET 8 = not_aux2
* NET 19 = mbk_buf_not_aux6
* NET 22 = not_y[2]
* NET 23 = not_aux6
* NET 26 = oa22_x2_3_sig
* NET 27 = z[4]
* NET 28 = o4_x2_sig
* NET 29 = not_y[0]
* NET 31 = o3_x2_sig
* NET 38 = mbk_buf_not_aux2
* NET 39 = not_aux9
* NET 40 = o2_x2_2_sig
* NET 54 = z[3]
* NET 59 = oa22_x2_2_sig
* NET 61 = nao2o22_x1_sig
* NET 64 = a4_x2_sig
* NET 67 = not_x[2]
* NET 68 = not_aux7
* NET 72 = not_aux3
* NET 74 = z[2]
* NET 82 = xr2_x1_2_sig
* NET 85 = not_x[0]
* NET 88 = o2_x2_sig
* NET 90 = not_aux4
* NET 91 = not_aux5
* NET 93 = no4_x1_sig
* NET 96 = no2_x1_sig
* NET 99 = aux2
* NET 105 = inv_x2_2_sig
* NET 109 = xr2_x1_4_sig
* NET 114 = mbk_buf_aux2
* NET 115 = xr2_x1_3_sig
* NET 124 = aux10
* NET 126 = nao22_x1_sig
* NET 129 = a3_x2_sig
* NET 131 = y[2]
* NET 135 = oa22_x2_sig
* NET 138 = inv_x2_sig
* NET 140 = vss
* NET 141 = z[0]
* NET 143 = z[1]
* NET 146 = aux0
* NET 149 = y[0]
* NET 151 = xr2_x1_sig
* NET 154 = aux1
* NET 156 = x[0]
* NET 158 = x[1]
* NET 161 = xr2_x1_5_sig
* NET 163 = x[2]
* NET 164 = y[1]
* NET 165 = a2_x2_sig
* NET 167 = vdd
Mtr_00314 153 158 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00313 167 154 155 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00312 151 153 152 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00311 152 154 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00310 152 155 151 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00309 167 158 152 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00308 154 157 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00307 167 156 157 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00306 157 164 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00305 165 166 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00304 167 164 166 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 166 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00302 159 158 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 167 165 160 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00300 161 159 162 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00299 162 165 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00298 162 160 161 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00297 167 158 162 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00296 167 148 143 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00295 144 151 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00294 147 149 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 145 149 148 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 148 147 144 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 167 154 145 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 141 142 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00289 167 146 142 167 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00288 146 150 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00287 167 149 150 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00286 150 156 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00285 138 158 167 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00284 167 161 134 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00283 129 134 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00282 167 126 134 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 134 135 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 167 133 135 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00279 104 131 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 104 138 133 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 133 164 104 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 124 120 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00275 167 156 120 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 120 131 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00273 106 124 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00272 167 114 108 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00271 109 106 101 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00270 101 114 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00269 101 108 109 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00268 167 124 101 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00267 105 124 167 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00266 113 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00265 167 114 119 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00264 115 113 102 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00263 102 114 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00262 102 119 115 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00261 167 163 102 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00260 167 124 126 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00259 103 164 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00258 126 163 103 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00257 167 91 95 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00256 94 96 92 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00255 92 149 93 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00254 95 90 94 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00253 87 129 89 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00252 167 93 87 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00251 88 89 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00250 99 100 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00249 167 158 100 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00248 100 164 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00247 97 164 96 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00246 167 131 97 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00245 84 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 167 131 86 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 82 84 83 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00242 83 131 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00241 83 86 82 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00240 167 163 83 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00239 77 78 79 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00238 167 75 80 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 76 149 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 79 109 76 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00235 80 115 77 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 81 82 80 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00233 79 85 81 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 74 79 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00231 78 85 167 167 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00230 167 149 75 167 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00229 85 156 167 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00228 114 98 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00227 167 99 98 167 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00226 50 72 66 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00225 167 67 50 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00224 68 66 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00223 91 69 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00222 167 85 69 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00221 69 131 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 52 158 71 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00219 167 164 52 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00218 72 71 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00217 90 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 167 72 90 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00215 167 53 54 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00214 43 88 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 43 59 53 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 53 149 43 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 64 62 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00210 62 85 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00209 167 131 62 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00208 62 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 167 158 62 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 167 57 59 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00205 45 64 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 45 61 57 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00203 57 156 45 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00202 42 39 41 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00201 167 156 42 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00200 40 41 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00199 167 163 39 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 39 38 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 39 131 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 33 29 32 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00195 34 67 33 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00194 30 91 34 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00193 167 38 30 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00192 167 32 28 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00191 67 163 167 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00190 167 149 35 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00189 35 39 36 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00188 36 85 37 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00187 31 37 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00186 61 68 25 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00185 25 22 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00184 24 131 61 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00183 167 23 24 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00182 167 40 27 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00181 27 28 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 167 26 27 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 27 31 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00178 167 21 26 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00177 20 105 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 20 68 21 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 21 19 20 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 167 99 8 167 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_00173 8 99 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00172 7 8 15 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00171 167 163 7 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00170 23 15 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00169 38 16 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00168 167 8 16 167 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00167 29 149 167 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00166 19 9 167 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00165 167 23 9 167 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00164 5 38 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00163 167 5 4 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00162 4 146 6 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00161 22 131 167 167 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00160 167 90 2 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00159 1 6 3 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00158 2 22 1 167 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00157 155 154 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00156 140 158 153 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00155 122 153 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 151 155 122 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00153 123 158 151 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 140 154 123 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 157 164 130 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 140 157 154 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 130 156 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00148 166 163 139 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 140 166 165 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 139 164 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00145 160 165 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00144 140 158 159 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00143 136 159 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 161 160 136 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 137 158 161 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 140 165 137 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 140 151 112 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00138 112 149 148 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00137 140 149 147 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00136 148 147 111 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00135 111 154 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00134 143 148 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00133 140 142 141 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00132 142 146 140 140 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00131 150 156 118 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00130 140 150 146 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 118 149 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 140 158 138 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00127 140 134 129 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 127 161 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 128 135 127 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 134 126 128 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00123 135 133 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00122 140 131 133 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00121 132 138 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00120 133 164 132 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00119 120 131 121 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 140 120 124 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 121 156 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 108 114 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00115 140 124 106 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00114 107 106 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 109 108 107 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 110 124 109 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 140 114 110 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 140 124 105 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 119 114 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00108 140 163 113 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 117 113 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 115 119 117 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 116 163 115 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 140 114 116 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 125 164 126 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 126 163 125 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 125 124 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 93 91 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00099 140 149 93 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00098 140 90 93 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00097 93 96 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00096 88 89 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 89 93 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00094 140 129 89 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00093 100 164 73 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00092 140 100 99 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 73 158 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 96 131 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00089 140 164 96 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00088 86 131 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00087 140 163 84 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00086 65 84 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 82 86 65 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00084 63 163 82 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 140 131 63 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 140 85 78 140 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00081 75 149 140 140 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00080 58 115 56 140 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00079 56 85 79 140 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00078 79 78 60 140 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00077 60 82 58 140 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00076 140 149 58 140 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00075 55 75 140 140 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00074 79 109 55 140 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00073 140 79 74 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 140 156 85 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 140 98 114 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 98 99 140 140 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00069 68 66 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 66 67 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00067 140 72 66 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00066 69 131 70 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 140 69 91 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 70 85 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 72 71 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 71 164 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00061 140 158 71 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00060 140 163 51 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 51 72 90 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 54 53 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 140 88 53 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 44 59 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00055 53 149 44 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 49 163 48 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 140 85 47 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 48 158 62 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 47 131 49 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 140 62 64 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 59 57 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 140 64 57 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 46 61 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 57 156 46 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 40 41 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 41 156 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00043 140 39 41 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00042 140 131 18 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 18 163 17 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 17 38 39 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 32 38 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 140 29 32 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00037 140 91 32 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00036 32 67 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00035 28 32 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 140 163 67 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 37 85 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 37 149 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00031 140 39 37 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00030 140 37 31 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 140 23 11 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 11 131 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 61 68 11 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 11 22 61 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 140 31 13 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 13 40 12 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 12 28 14 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 14 26 27 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 26 21 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 140 105 21 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00019 10 68 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 21 19 10 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 140 99 8 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 8 99 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 23 15 140 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 15 163 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 140 8 15 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 140 16 38 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 16 8 140 140 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00010 140 149 29 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 140 9 19 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 9 23 140 140 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00007 140 38 5 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 6 5 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 140 146 6 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 140 131 22 140 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 140 22 3 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 3 90 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 3 6 140 140 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C170 3 140 4.843e-14
C168 5 140 1.677e-14
C167 6 140 5.428e-14
C164 8 140 8.098e-14
C163 9 140 1.568e-14
C161 11 140 7.43e-15
C157 15 140 1.8635e-14
C156 16 140 1.568e-14
C152 19 140 4.839e-14
C151 20 140 6.05e-15
C150 21 140 1.767e-14
C149 22 140 7.915e-14
C148 23 140 1.2419e-13
C145 26 140 6.572e-14
C144 27 140 4.427e-14
C143 28 140 6.004e-14
C142 29 140 5.139e-14
C140 31 140 6.452e-14
C139 32 140 2.72e-14
C134 37 140 2.455e-14
C133 38 140 1.3676e-13
C132 39 140 8.026e-14
C131 40 140 8.126e-14
C130 41 140 1.8635e-14
C128 43 140 6.05e-15
C126 45 140 6.05e-15
C117 53 140 1.767e-14
C116 54 140 3.023e-14
C113 57 140 1.767e-14
C112 58 140 7.56e-15
C111 59 140 4.877e-14
C109 61 140 5.537e-14
C108 62 140 2.306e-14
C106 64 140 5.981e-14
C104 66 140 1.8635e-14
C103 67 140 8.878e-14
C102 68 140 9.75e-14
C101 69 140 1.8635e-14
C99 71 140 1.8635e-14
C98 72 140 8.447e-14
C95 74 140 2.469e-14
C94 75 140 2.378e-14
C91 78 140 2.128e-14
C90 79 140 3.608e-14
C89 80 140 7.56e-15
C87 82 140 4.51e-14
C86 83 140 9.7e-15
C85 84 140 2.596e-14
C84 85 140 1.796e-13
C83 86 140 2.16e-14
C81 88 140 8.305e-14
C80 89 140 1.8635e-14
C79 90 140 1.3453e-13
C78 91 140 1.0079e-13
C76 93 140 6.397e-14
C73 96 140 5.176e-14
C71 98 140 1.568e-14
C70 99 140 1.2586e-13
C69 100 140 1.8635e-14
C68 101 140 9.7e-15
C67 102 140 9.7e-15
C65 104 140 6.05e-15
C63 105 140 8.045e-14
C62 106 140 2.596e-14
C60 108 140 2.16e-14
C59 109 140 5.856e-14
C55 113 140 2.596e-14
C54 114 140 1.3106e-13
C53 115 140 5.966e-14
C49 119 140 2.16e-14
C48 120 140 1.8635e-14
C44 124 140 1.3855e-13
C43 125 140 4.11e-15
C42 126 140 5.027e-14
C39 129 140 5.925e-14
C37 131 140 3.5532e-13
C35 133 140 1.767e-14
C34 134 140 2.605e-14
C33 135 140 4.817e-14
C30 138 140 4.569e-14
C28 140 140 1.81812e-12
C27 141 140 2.371e-14
C26 142 140 1.568e-14
C25 143 140 3.815e-14
C22 146 140 1.5981e-13
C21 147 140 2.356e-14
C20 148 140 1.932e-14
C19 149 140 3.3457e-13
C18 150 140 1.8635e-14
C17 151 140 6.891e-14
C16 152 140 9.7e-15
C15 153 140 2.596e-14
C14 154 140 9.561e-14
C13 155 140 2.16e-14
C12 156 140 2.8771e-13
C11 157 140 1.8635e-14
C10 158 140 2.7737e-13
C9 159 140 2.596e-14
C8 160 140 2.16e-14
C7 161 140 5.485e-14
C6 162 140 9.7e-15
C5 163 140 4.0784e-13
C4 164 140 2.9152e-13
C3 165 140 5.409e-14
C2 166 140 1.8635e-14
C1 167 140 1.91192e-12
.ends mul3b_cougar

