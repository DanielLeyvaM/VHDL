* Spice description of act4_cougar
* Spice driver version -1209221468
* Date ( dd/mm/yyyy hh:mm:ss ): 22/11/2020 at 11:09:04

* INTERF clk dh[0] dh[1] dh[2] dh[3] dm[0] dm[1] dm[2] dm[3] rst uh[0] uh[1] 
* INTERF uh[2] uh[3] um[0] um[1] um[2] um[3] vdd vss 


.subckt act4_cougar 604 180 124 17 74 408 363 324 260 595 225 224 228 182 563 499 588 497 608 561 
* NET 17 = dh[2]
* NET 18 = mdh_2_ins.ckr
* NET 19 = mdh_2_ins.nckr
* NET 20 = mdh_2_ins.sff_m
* NET 21 = mdh_2_ins.y
* NET 23 = mdh_2_ins.sff_s
* NET 25 = mdh_2_ins.u
* NET 28 = no2_x1_sig
* NET 32 = nxr2_x1_sig
* NET 35 = mdm_1_ins.ckr
* NET 36 = mdm_1_ins.nckr
* NET 37 = mdm_1_ins.sff_m
* NET 39 = mdm_1_ins.sff_s
* NET 42 = mdm_1_ins.y
* NET 45 = mdm_1_ins.u
* NET 50 = mdm_3_ins.ckr
* NET 51 = mdm_3_ins.nckr
* NET 52 = mdm_3_ins.sff_s
* NET 54 = mdm_3_ins.sff_m
* NET 55 = mdm_3_ins.y
* NET 60 = mdm_3_ins.u
* NET 62 = no2_x1_8_sig
* NET 64 = na2_x1_4_sig
* NET 66 = noa22_x1_5_sig
* NET 71 = o3_x2_2_sig
* NET 74 = dh[3]
* NET 76 = mdh[2]
* NET 79 = mbk_buf_aux14
* NET 80 = no2_x1_4_sig
* NET 84 = no4_x1_2_sig
* NET 85 = noa2a2a23_x1_sig
* NET 86 = muh_1_ins.y
* NET 88 = muh_1_ins.sff_s
* NET 90 = no2_x1_3_sig
* NET 91 = muh_1_ins.u
* NET 92 = muh_1_ins.sff_m
* NET 94 = muh_1_ins.ckr
* NET 95 = muh_1_ins.nckr
* NET 98 = nxr2_x1_4_sig
* NET 102 = not_aux35
* NET 103 = no3_x1_2_sig
* NET 104 = mbk_buf_mdm[3]
* NET 105 = no2_x1_7_sig
* NET 124 = dh[1]
* NET 128 = not_mdh[2]
* NET 130 = an12_x1_sig
* NET 135 = nxr2_x1_2_sig
* NET 136 = mdh[3]
* NET 138 = mdh_3_ins.sff_s
* NET 139 = mdh_3_ins.y
* NET 141 = no2_x1_2_sig
* NET 142 = mdh_3_ins.u
* NET 143 = mdh_3_ins.sff_m
* NET 145 = mdh_3_ins.ckr
* NET 147 = mdh_3_ins.nckr
* NET 148 = nao22_x1_sig
* NET 151 = a3_x2_2_sig
* NET 153 = inv_x2_2_sig
* NET 155 = aux23
* NET 157 = mdm_2_ins.y
* NET 159 = mdm_2_ins.sff_s
* NET 160 = mdm_2_ins.ckr
* NET 161 = mdm_2_ins.u
* NET 164 = mdm_2_ins.sff_m
* NET 166 = mdm_2_ins.nckr
* NET 169 = noa22_x1_6_sig
* NET 172 = on12_x1_6_sig
* NET 173 = xr2_x1_6_sig
* NET 180 = dh[0]
* NET 182 = uh[3]
* NET 183 = aux14
* NET 184 = not_aux11
* NET 185 = not_muh[3]
* NET 188 = na2_x1_3_sig
* NET 190 = no3_x1_sig
* NET 192 = o2_x2_3_sig
* NET 195 = not_boom_init_9
* NET 198 = muh_0_ins.sff_s
* NET 200 = muh_0_ins.y
* NET 202 = muh_0_ins.sff_m
* NET 204 = muh_0_ins.u
* NET 205 = muh_0_ins.ckr
* NET 206 = muh_0_ins.nckr
* NET 208 = mbk_buf_not_aux22
* NET 210 = o2_x2_4_sig
* NET 224 = uh[1]
* NET 225 = uh[0]
* NET 228 = uh[2]
* NET 232 = a2_x2_2_sig
* NET 233 = muh[1]
* NET 235 = muh_3_ins.y
* NET 236 = muh_3_ins.sff_m
* NET 239 = muh_3_ins.sff_s
* NET 240 = muh_3_ins.u
* NET 242 = muh_3_ins.ckr
* NET 243 = muh_3_ins.nckr
* NET 245 = on12_x1_4_sig
* NET 246 = noa22_x1_3_sig
* NET 248 = na2_x1_2_sig
* NET 250 = not_aux18
* NET 251 = mdm[1]
* NET 252 = not_mdm[2]
* NET 256 = no4_x1_sig
* NET 258 = aux35
* NET 260 = dm[3]
* NET 261 = inv_x2_sig
* NET 268 = a3_x2_sig
* NET 271 = not_aux24
* NET 276 = noa22_x1_4_sig
* NET 283 = xr2_x1_5_sig
* NET 286 = na4_x1_2_sig
* NET 289 = not_aux22
* NET 296 = xr2_x1_3_sig
* NET 297 = not_mdm[1]
* NET 305 = not_muh[1]
* NET 307 = on12_x1_5_sig
* NET 308 = na3_x1_2_sig
* NET 314 = muh[3]
* NET 315 = no2_x1_5_sig
* NET 322 = mbk_buf_not_aux19
* NET 323 = muh[0]
* NET 324 = dm[2]
* NET 326 = na3_x1_sig
* NET 329 = na2_x1_sig
* NET 330 = mdm[2]
* NET 331 = na4_x1_sig
* NET 332 = not_muh[2]
* NET 335 = xr2_x1_4_sig
* NET 338 = muh[2]
* NET 340 = muh_2_ins.sff_s
* NET 341 = muh_2_ins.y
* NET 343 = muh_2_ins.sff_m
* NET 344 = ao22_x2_sig
* NET 345 = muh_2_ins.u
* NET 347 = muh_2_ins.ckr
* NET 348 = muh_2_ins.nckr
* NET 349 = aux26
* NET 352 = an12_x1_3_sig
* NET 353 = mbk_buf_not_aux1
* NET 354 = not_aux1
* NET 357 = not_aux19
* NET 358 = not_aux38
* NET 361 = not_mdm[0]
* NET 362 = aux40
* NET 363 = dm[1]
* NET 371 = no4_x1_3_sig
* NET 376 = aux1
* NET 384 = not_aux9
* NET 388 = inv_x2_3_sig
* NET 390 = not_aux31
* NET 395 = a4_x2_sig
* NET 396 = an12_x1_2_sig
* NET 397 = a2_x2_sig
* NET 400 = not_mdh[1]
* NET 404 = aux37
* NET 407 = mbk_buf_not_aux9
* NET 408 = dm[0]
* NET 412 = mdm[3]
* NET 413 = mdm_0_ins.sff_s
* NET 415 = mdm_0_ins.ckr
* NET 416 = mdm_0_ins.sff_m
* NET 418 = mdm_0_ins.y
* NET 419 = mdm_0_ins.u
* NET 420 = no2_x1_6_sig
* NET 421 = mdm_0_ins.nckr
* NET 425 = mdm[0]
* NET 426 = nxr2_x1_3_sig
* NET 429 = aux10
* NET 432 = mbk_buf_aux10
* NET 435 = mdh[1]
* NET 436 = mdh_1_ins.sff_s
* NET 438 = mdh_1_ins.y
* NET 440 = mdh_1_ins.sff_m
* NET 442 = xr2_x1_2_sig
* NET 443 = mdh_1_ins.u
* NET 444 = mdh_1_ins.ckr
* NET 445 = mdh_1_ins.nckr
* NET 447 = on12_x1_3_sig
* NET 448 = o2_x2_2_sig
* NET 449 = o3_x2_sig
* NET 450 = noa22_x1_2_sig
* NET 451 = on12_x1_2_sig
* NET 455 = mum_1_ins.sff_s
* NET 456 = mum_1_ins.y
* NET 458 = mum_1_ins.sff_m
* NET 459 = mum_1_ins.u
* NET 461 = mum_1_ins.ckr
* NET 462 = mum[1]
* NET 463 = mum_1_ins.nckr
* NET 466 = not_aux25
* NET 470 = o3_x2_3_sig
* NET 471 = noa22_x1_7_sig
* NET 473 = o2_x2_5_sig
* NET 479 = not_mum[1]
* NET 483 = aux34
* NET 497 = um[3]
* NET 499 = um[1]
* NET 502 = mum_3_ins.y
* NET 503 = mum_3_ins.sff_s
* NET 505 = mum_3_ins.u
* NET 507 = mum_3_ins.sff_m
* NET 510 = mum_3_ins.ckr
* NET 511 = mum_3_ins.nckr
* NET 513 = not_aux0
* NET 514 = not_mdh[0]
* NET 517 = mum[3]
* NET 521 = xr2_x1_8_sig
* NET 527 = noa22_x1_9_sig
* NET 530 = not_mum[3]
* NET 532 = o2_x2_7_sig
* NET 533 = o3_x2_4_sig
* NET 534 = on12_x1_8_sig
* NET 537 = oa22_x2_sig
* NET 538 = mbk_buf_mum[1]
* NET 542 = xr2_x1_7_sig
* NET 546 = on12_x1_7_sig
* NET 551 = mum_2_ins.sff_m
* NET 552 = mum_2_ins.sff_s
* NET 553 = mum_2_ins.y
* NET 555 = noa22_x1_8_sig
* NET 557 = mum_2_ins.u
* NET 558 = mum_2_ins.ckr
* NET 559 = mum_2_ins.nckr
* NET 561 = vss
* NET 563 = um[0]
* NET 564 = aux9
* NET 567 = mbk_buf_aux9
* NET 570 = xr2_x1_sig
* NET 571 = aux0
* NET 573 = o2_x2_sig
* NET 574 = on12_x1_sig
* NET 577 = mdh[0]
* NET 578 = mdh_0_ins.sff_s
* NET 579 = mdh_0_ins.y
* NET 581 = mdh_0_ins.sff_m
* NET 582 = noa22_x1_sig
* NET 583 = mdh_0_ins.u
* NET 585 = mdh_0_ins.ckr
* NET 586 = mdh_0_ins.nckr
* NET 588 = um[2]
* NET 589 = not_mum[0]
* NET 592 = o2_x2_6_sig
* NET 593 = mum[2]
* NET 594 = not_mum[2]
* NET 595 = rst
* NET 598 = mum[0]
* NET 599 = mum_0_ins.sff_s
* NET 600 = mum_0_ins.y
* NET 602 = mum_0_ins.sff_m
* NET 603 = no2_x1_9_sig
* NET 604 = clk
* NET 606 = mum_0_ins.u
* NET 607 = mum_0_ins.ckr
* NET 608 = vdd
* NET 609 = mum_0_ins.nckr
Mtr_01214 597 598 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01213 599 607 597 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01212 600 609 599 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01211 602 609 601 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01210 601 600 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01209 605 607 602 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01208 609 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01207 608 609 607 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01206 606 603 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01205 608 606 605 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01204 608 599 598 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01203 598 599 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01202 600 602 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01201 591 594 590 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01200 608 598 591 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01199 592 590 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01198 596 598 603 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01197 608 595 596 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01196 566 577 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01195 608 567 568 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01194 570 566 569 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01193 569 567 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01192 569 568 570 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01191 608 577 569 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01190 567 565 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01189 608 564 565 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01188 594 593 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01187 588 587 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01186 608 593 587 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01185 589 598 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01184 608 595 575 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01183 582 574 575 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01182 575 573 582 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01181 576 577 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01180 578 585 576 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01179 579 586 578 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01178 581 586 580 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01177 580 579 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01176 584 585 581 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01175 586 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01174 608 586 585 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01173 583 582 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01172 608 583 584 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01171 608 578 577 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01170 577 578 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01169 579 581 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01168 563 562 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01167 608 598 562 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01166 608 570 574 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01165 574 572 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01164 608 571 572 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01163 518 517 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01162 608 538 524 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01161 521 518 488 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01160 488 538 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01159 488 524 521 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01158 608 517 488 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01157 608 542 546 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01156 546 543 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01155 608 589 543 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01154 494 593 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01153 552 558 494 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01152 553 559 552 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01151 551 559 495 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01150 495 553 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01149 496 558 551 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01148 559 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01147 608 559 558 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01146 557 555 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01145 608 557 496 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01144 608 552 593 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01143 593 552 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01142 553 551 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01141 540 538 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01140 608 593 545 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01139 542 540 492 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01138 492 593 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01137 492 545 542 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01136 608 538 492 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01135 608 595 493 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01134 555 546 493 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01133 493 592 555 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01132 490 530 531 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01131 608 598 490 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01130 532 531 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01129 499 500 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01128 608 538 500 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01127 608 521 534 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01126 534 522 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01125 608 594 522 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01124 608 595 489 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01123 527 537 489 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01122 489 532 527 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01121 608 536 537 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01120 491 589 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01119 491 533 536 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01118 536 534 491 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01117 513 571 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01116 497 498 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01115 608 517 498 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01114 484 517 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01113 503 510 484 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01112 502 511 503 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01111 507 511 486 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01110 486 502 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01109 485 510 507 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01108 511 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01107 608 511 510 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01106 505 527 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01105 608 505 485 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01104 608 503 517 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01103 517 503 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01102 502 507 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01101 487 514 515 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01100 608 513 487 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01099 573 515 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01098 514 577 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01097 608 593 480 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01096 481 538 482 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01095 482 530 483 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01094 480 589 481 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01093 608 530 476 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01092 476 593 477 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01091 477 479 478 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01090 533 478 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01089 538 464 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01088 608 462 464 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01087 479 538 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01086 474 479 475 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01085 608 598 474 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01084 473 475 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01083 466 465 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01082 608 594 465 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01081 465 517 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01080 608 595 472 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01079 471 470 472 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01078 472 473 471 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01077 608 466 467 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01076 467 538 469 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01075 469 589 468 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01074 470 468 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01073 608 449 451 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01072 451 453 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01071 608 595 453 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01070 454 462 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01069 455 461 454 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01068 456 463 455 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01067 458 463 457 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01066 457 456 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01065 460 461 458 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01064 463 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01063 608 463 461 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01062 459 471 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01061 608 459 460 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01060 608 455 462 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01059 462 455 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01058 456 458 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01057 437 435 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01056 436 444 437 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01055 438 445 436 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01054 440 445 439 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01053 439 438 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01052 441 444 440 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01051 445 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01050 608 445 444 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01049 443 450 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01048 608 443 441 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01047 608 436 435 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01046 435 436 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01045 438 440 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01044 432 430 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01043 608 429 430 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01042 608 451 452 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01041 450 447 452 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01040 452 448 450 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01039 431 435 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01038 608 432 433 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01037 442 431 434 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01036 434 432 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01035 434 433 442 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01034 608 435 434 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01033 608 442 447 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01032 447 446 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01031 608 571 446 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01030 608 423 383 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01029 383 424 426 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01028 383 483 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01027 426 425 383 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01026 608 483 424 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01025 423 425 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01024 378 425 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01023 413 415 378 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01022 418 421 413 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01021 416 421 377 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01020 377 418 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01019 380 415 416 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01018 421 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01017 608 421 415 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01016 419 420 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01015 608 419 380 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01014 608 413 425 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01013 425 413 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01012 418 416 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01011 530 517 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01010 382 426 420 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01009 608 595 382 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01008 375 462 376 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01007 608 412 375 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01006 408 405 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01005 608 425 405 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01004 372 400 398 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01003 608 513 372 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01002 448 398 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01001 608 577 373 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01000 373 407 374 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00999 374 404 401 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00998 449 401 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00997 384 564 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00996 407 406 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00995 608 384 406 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00994 395 385 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00993 385 514 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00992 608 435 385 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00991 385 390 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00990 608 388 385 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00989 397 391 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00988 608 390 391 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00987 391 513 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00986 364 384 429 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00985 608 514 364 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00984 388 404 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00983 608 397 368 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00982 370 396 369 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00981 369 595 371 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00980 368 395 370 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00979 351 362 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00978 608 351 350 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00977 350 353 352 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00976 355 354 357 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00975 608 530 355 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00974 354 376 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00973 608 358 360 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00972 359 589 362 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00971 360 361 359 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00970 353 356 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00969 608 354 356 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00968 361 425 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00967 608 466 349 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00966 349 362 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00965 349 376 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00964 608 332 331 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00963 331 330 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00962 608 376 331 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00961 331 425 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00960 339 338 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00959 340 347 339 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00958 341 348 340 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00957 343 348 342 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00956 342 341 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00955 346 347 343 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00954 348 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00953 608 348 347 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00952 345 344 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00951 608 345 346 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00950 608 340 338 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00949 338 340 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00948 341 343 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00947 608 336 344 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00946 336 371 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00945 608 335 337 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00944 337 349 336 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00943 608 338 332 608 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_00942 332 338 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00941 324 325 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00940 608 330 325 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00939 329 598 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00938 608 594 329 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00937 608 326 328 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00936 327 331 564 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00935 328 329 327 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00934 334 349 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00933 608 334 333 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00932 333 338 396 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00931 320 322 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00930 608 323 321 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00929 296 320 293 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00928 293 323 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00927 293 321 296 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00926 608 322 293 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00925 608 338 286 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00924 286 517 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00923 608 352 286 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00922 286 323 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00921 289 318 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00920 318 357 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00919 608 598 318 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00918 318 594 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00917 608 425 318 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00916 284 286 315 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00915 608 593 284 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00914 322 319 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00913 608 357 319 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00912 311 314 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00911 608 315 312 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00910 283 311 281 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00909 281 315 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00908 281 312 283 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00907 608 314 281 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00906 608 283 307 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00905 307 279 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00904 608 305 279 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00903 608 595 275 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00902 276 307 275 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00901 275 308 276 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00900 608 330 300 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00899 268 300 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00898 608 271 300 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00897 300 425 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00896 608 407 308 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00895 308 305 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00894 308 314 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00893 608 517 326 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00892 326 297 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00891 326 323 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00890 271 304 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00889 608 332 304 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00888 304 323 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00887 261 429 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00886 571 314 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00885 608 305 571 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00884 390 298 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00883 298 268 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00882 608 297 298 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00881 298 594 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00880 608 598 298 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00879 257 483 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00878 608 257 259 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00877 259 361 258 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00876 248 250 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00875 608 296 248 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00874 608 361 253 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00873 254 251 255 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00872 255 252 256 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00871 253 593 254 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00870 608 595 247 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00869 246 248 247 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00868 247 245 246 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00867 250 249 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00866 608 598 249 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00865 249 256 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00864 608 323 245 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00863 245 244 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00862 608 250 244 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00861 231 338 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00860 608 232 234 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00859 335 231 230 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00858 230 232 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00857 230 234 335 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00856 608 338 230 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00855 238 314 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00854 239 242 238 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00853 235 243 239 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00852 236 243 237 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00851 237 235 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00850 241 242 236 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00849 243 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00848 608 243 242 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00847 240 276 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00846 608 240 241 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00845 608 239 314 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00844 314 239 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00843 235 236 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00842 305 233 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00841 232 229 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00840 608 323 229 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00839 229 233 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00838 400 435 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00837 225 222 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00836 608 323 222 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00835 228 227 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00834 608 338 227 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00833 363 226 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00832 608 251 226 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00831 224 223 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00830 608 233 223 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00829 208 207 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00828 608 289 207 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00827 165 323 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00826 198 205 165 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00825 200 206 198 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00824 202 206 167 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00823 167 200 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00822 168 205 202 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00821 206 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00820 608 206 205 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00819 204 246 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00818 608 204 168 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00817 608 198 323 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00816 323 198 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00815 200 202 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00814 176 208 209 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00813 608 358 176 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00812 210 209 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00811 178 252 211 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00810 608 251 178 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00809 358 211 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00808 297 251 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00807 608 314 149 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00806 150 577 190 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00805 149 400 150 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00804 608 233 404 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00803 404 185 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00802 404 184 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00801 152 195 191 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00800 608 271 152 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00799 192 191 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00798 608 193 156 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00797 156 194 195 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00796 156 323 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00795 195 233 156 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00794 608 323 194 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00793 193 233 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00792 188 271 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00791 608 314 188 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00790 180 179 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00789 608 577 179 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00788 185 314 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00787 182 181 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00786 608 314 181 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00785 608 233 132 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00784 134 400 133 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00783 133 261 183 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00782 132 185 134 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00781 252 330 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00780 608 595 170 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00779 169 172 170 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00778 170 210 169 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00777 155 330 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00776 608 289 155 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00775 608 173 172 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00774 172 171 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00773 608 297 171 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00772 175 330 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00771 608 258 177 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00770 173 175 174 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00769 174 258 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00768 174 177 173 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00767 608 330 174 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00766 153 155 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00765 608 153 154 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00764 151 154 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00763 608 192 154 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00762 154 297 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00761 158 330 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00760 159 160 158 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00759 157 166 159 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00758 164 166 162 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00757 162 157 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00756 163 160 164 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00755 166 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00754 608 166 160 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00753 161 169 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00752 608 161 163 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00751 608 159 330 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00750 330 159 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00749 157 164 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00748 608 151 148 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00747 146 190 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00746 148 195 146 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00745 608 123 126 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00744 126 125 135 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00743 126 130 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00742 135 136 126 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00741 608 130 125 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00740 123 136 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00739 131 135 141 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00738 608 595 131 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00737 127 183 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00736 608 127 129 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00735 129 128 130 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00734 137 136 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00733 138 145 137 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00732 139 147 138 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00731 143 147 140 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00730 140 139 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00729 144 145 143 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00728 147 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00727 608 147 145 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00726 142 141 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00725 608 142 144 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00724 608 138 136 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00723 136 138 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00722 139 143 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00721 124 122 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00720 608 435 122 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00719 608 102 68 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00718 69 297 103 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00717 68 252 69 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00716 72 252 105 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00715 608 104 72 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00714 608 97 67 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00713 67 100 98 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00712 67 103 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00711 98 104 67 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00710 608 103 100 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00709 97 104 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00708 104 96 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00707 608 412 96 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00706 59 233 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00705 88 94 59 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00704 86 95 88 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00703 92 95 58 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00702 58 86 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00701 61 94 92 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00700 95 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00699 608 95 94 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00698 91 90 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00697 608 91 61 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00696 608 88 233 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00695 233 88 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00694 86 92 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00693 49 85 90 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00692 608 595 49 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00691 260 73 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00690 608 104 73 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00689 608 233 48 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00688 47 195 46 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00687 46 155 84 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00686 48 251 47 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00685 41 148 85 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00684 85 233 41 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00683 41 188 40 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00682 40 84 41 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00681 608 233 40 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00680 40 80 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00679 34 195 80 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00678 608 184 34 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00677 128 76 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00676 608 183 78 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00675 608 78 79 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00674 79 78 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00673 77 128 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00672 608 77 27 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00671 27 136 184 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00670 74 75 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00669 608 136 75 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00668 608 102 15 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00667 15 251 14 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00666 14 105 70 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00665 71 70 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00664 53 412 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00663 52 50 53 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00662 55 51 52 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00661 54 51 56 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00660 56 55 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00659 57 50 54 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00658 51 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00657 608 51 50 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00656 60 62 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00655 608 60 57 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00654 608 52 412 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00653 412 52 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00652 55 54 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00651 63 98 62 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00650 608 595 63 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00649 608 595 65 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00648 66 71 65 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00647 65 64 66 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00646 102 258 608 608 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00645 64 102 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00644 608 251 64 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00643 38 251 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00642 39 35 38 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00641 42 36 39 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00640 37 36 44 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00639 44 42 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00638 43 35 37 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00637 36 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00636 608 36 35 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00635 45 66 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00634 608 45 43 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00633 608 39 251 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00632 251 39 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00631 42 37 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00630 608 30 33 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00629 33 31 32 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00628 33 79 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00627 32 76 33 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00626 608 79 31 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00625 30 76 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00624 17 16 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00623 608 76 16 608 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00622 29 32 28 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00621 608 595 29 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00620 24 76 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00619 23 18 24 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00618 21 19 23 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00617 20 19 22 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00616 22 21 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00615 26 18 20 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00614 19 604 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00613 608 19 18 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00612 25 28 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00611 608 25 26 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00610 608 23 76 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00609 76 23 608 608 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00608 21 20 608 608 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00607 549 609 599 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00606 561 598 549 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00605 599 607 600 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00604 561 600 554 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00603 554 607 602 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00602 602 609 560 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00601 607 609 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00600 561 604 609 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00599 560 606 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00598 561 603 606 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00597 598 599 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00596 561 599 598 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00595 600 602 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00594 592 590 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00593 590 598 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00592 561 594 590 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00591 603 595 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00590 561 598 603 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00589 568 567 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00588 561 577 566 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00587 504 566 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00586 570 568 504 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00585 509 577 570 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00584 561 567 509 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00583 561 565 567 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00582 565 564 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00581 561 593 594 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00580 561 587 588 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00579 587 593 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00578 561 598 589 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00577 561 574 516 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00576 516 573 582 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00575 582 595 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00574 520 586 578 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00573 561 577 520 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00572 578 585 579 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00571 561 579 526 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00570 526 585 581 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00569 581 586 529 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00568 585 586 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00567 561 604 586 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00566 529 583 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00565 561 582 583 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00564 577 578 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00563 561 578 577 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00562 579 581 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00561 561 562 563 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00560 562 598 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00559 572 571 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00558 512 570 574 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00557 561 572 512 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00556 524 538 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00555 561 517 518 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00554 519 518 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00553 521 524 519 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00552 525 517 521 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00551 561 538 525 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00550 543 589 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00549 544 542 546 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00548 561 543 544 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00547 548 559 552 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00546 561 593 548 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00545 552 558 553 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00544 561 553 550 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00543 550 558 551 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00542 551 559 556 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00541 558 559 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00540 561 604 559 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00539 556 557 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00538 561 555 557 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00537 593 552 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00536 561 552 593 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00535 553 551 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00534 545 593 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00533 561 538 540 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00532 541 540 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00531 542 545 541 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00530 539 538 542 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00529 561 593 539 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00528 561 546 547 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00527 547 592 555 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00526 555 595 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00525 532 531 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00524 531 598 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00523 561 530 531 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00522 561 500 499 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00521 500 538 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00520 522 594 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00519 523 521 534 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00518 561 522 523 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00517 561 537 528 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00516 528 532 527 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00515 527 595 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00514 537 536 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00513 561 589 536 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00512 535 533 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00511 536 534 535 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00510 561 571 513 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00509 561 498 497 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00508 498 517 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00507 501 511 503 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00506 561 517 501 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00505 503 510 502 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00504 561 502 506 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00503 506 510 507 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00502 507 511 508 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00501 510 511 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00500 561 604 511 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00499 508 505 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00498 561 527 505 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00497 517 503 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00496 561 503 517 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00495 502 507 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00494 573 515 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00493 515 513 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00492 561 514 515 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00491 561 577 514 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00490 483 593 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00489 561 530 483 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00488 561 589 483 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00487 483 538 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00486 478 479 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00485 478 530 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00484 561 593 478 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00483 561 478 533 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00482 561 464 538 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00481 464 462 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00480 561 538 479 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00479 473 475 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00478 475 598 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00477 561 479 475 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00476 465 517 414 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00475 561 465 466 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00474 414 594 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00473 561 470 422 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00472 422 473 471 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00471 471 595 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00470 468 589 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00469 468 466 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00468 561 538 468 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00467 561 468 470 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00466 453 595 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00465 402 449 451 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00464 561 453 402 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00463 410 463 455 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00462 561 462 410 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00461 455 461 456 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00460 561 456 409 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00459 409 461 458 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00458 458 463 411 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00457 461 463 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00456 561 604 463 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00455 411 459 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00454 561 471 459 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00453 462 455 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00452 561 455 462 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00451 456 458 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00450 389 445 436 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00449 561 435 389 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00448 436 444 438 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00447 561 438 393 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00446 393 444 440 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00445 440 445 394 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00444 444 445 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00443 561 604 445 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00442 394 443 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00441 561 450 443 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00440 435 436 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00439 561 436 435 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00438 438 440 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00437 561 430 432 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00436 430 429 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00435 561 447 403 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00434 403 448 450 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00433 450 451 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00432 433 432 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00431 561 435 431 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00430 386 431 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00429 442 433 386 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00428 387 435 442 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00427 561 432 387 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00426 446 571 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00425 399 442 447 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00424 561 446 399 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00423 561 483 428 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00422 428 423 426 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00421 426 424 427 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00420 427 425 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00419 561 425 423 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00418 424 483 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00417 379 421 413 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00416 561 425 379 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00415 413 415 418 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00414 561 418 417 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00413 417 415 416 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00412 416 421 381 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00411 415 421 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00410 561 604 421 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00409 381 419 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00408 561 420 419 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00407 425 413 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00406 561 413 425 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00405 418 416 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00404 561 517 530 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00403 420 595 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00402 561 426 420 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00401 376 412 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00400 561 462 376 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00399 561 405 408 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00398 405 425 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00397 448 398 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00396 398 513 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00395 561 400 398 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00394 401 404 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00393 401 577 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00392 561 407 401 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00391 561 401 449 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00390 561 564 384 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00389 561 406 407 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00388 406 384 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00387 365 390 367 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00386 561 514 366 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00385 367 388 385 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 366 435 365 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00383 561 385 395 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 391 513 392 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 561 391 397 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 392 390 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00379 429 514 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00378 561 384 429 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00377 561 404 388 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00376 371 397 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00375 561 595 371 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00374 561 395 371 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00373 371 396 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00372 561 362 351 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00371 352 351 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00370 561 353 352 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00369 357 530 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00368 561 354 357 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00367 561 376 354 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00366 561 361 362 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00365 362 358 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00364 362 589 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00363 561 356 353 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00362 356 354 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00361 561 425 361 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00360 561 376 317 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00359 317 466 316 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00358 316 362 349 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00357 561 425 303 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00356 303 332 302 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00355 302 330 301 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00354 301 376 331 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00353 309 348 340 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00352 561 338 309 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00351 340 347 341 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00350 561 341 310 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00349 310 347 343 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00348 343 348 313 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00347 347 348 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00346 561 604 348 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00345 313 345 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00344 561 344 345 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00343 338 340 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00342 561 340 338 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00341 341 343 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00340 336 335 306 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00339 306 349 336 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00338 561 371 306 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00337 344 336 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00336 561 338 332 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00335 332 338 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 561 325 324 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00333 325 330 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00332 561 598 299 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00331 299 594 329 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00330 561 329 564 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00329 564 326 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00328 564 331 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00327 561 349 334 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00326 396 334 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00325 561 338 396 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00324 321 323 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00323 561 322 320 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00322 295 320 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00321 296 321 295 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00320 294 322 296 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00319 561 323 294 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00318 561 323 288 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00317 288 338 287 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00316 287 517 285 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00315 285 352 286 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00314 291 594 290 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00313 561 357 292 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00312 290 425 318 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00311 292 598 291 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00310 561 318 289 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00309 315 593 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00308 561 286 315 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00307 561 319 322 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00306 319 357 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00305 312 315 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00304 561 314 311 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00303 280 311 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00302 283 312 280 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 282 314 283 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00300 561 315 282 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00299 279 305 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00298 278 283 307 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00297 561 279 278 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00296 561 307 277 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 277 308 276 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00294 276 595 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 561 300 268 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 269 330 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 267 425 269 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 300 271 267 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 561 314 274 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00288 274 407 273 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00287 273 305 308 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00286 561 323 263 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00285 263 517 262 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00284 262 297 326 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00283 304 323 270 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00282 561 304 271 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 270 332 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 561 429 261 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00279 561 314 272 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 272 305 571 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 264 594 266 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 561 268 265 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 266 598 298 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 265 297 264 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00273 561 298 390 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00272 561 483 257 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00271 258 257 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00270 561 361 258 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00269 561 250 220 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 220 296 248 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 256 361 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00266 561 252 256 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00265 561 593 256 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00264 256 251 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00263 561 248 219 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 219 245 246 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 246 595 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 249 256 221 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00259 561 249 250 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00258 221 598 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00257 244 250 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00256 218 323 245 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00255 561 244 218 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00254 234 232 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00253 561 338 231 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00252 213 231 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00251 335 234 213 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00250 214 338 335 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00249 561 232 214 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00248 215 243 239 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00247 561 314 215 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00246 239 242 235 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00245 561 235 216 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00244 216 242 236 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00243 236 243 217 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00242 242 243 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00241 561 604 243 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00240 217 240 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00239 561 276 240 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00238 314 239 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 561 239 314 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 235 236 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00235 561 233 305 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 229 233 212 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00233 561 229 232 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 212 323 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 561 435 400 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 561 222 225 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 222 323 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00228 561 227 228 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00227 227 338 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00226 561 226 363 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00225 226 251 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00224 561 223 224 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00223 223 233 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00222 561 207 208 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00221 207 289 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00220 199 206 198 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00219 561 323 199 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00218 198 205 200 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00217 561 200 201 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00216 201 205 202 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00215 202 206 203 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00214 205 206 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00213 561 604 206 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00212 203 204 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00211 561 246 204 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00210 323 198 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00209 561 198 323 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00208 200 202 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00207 210 209 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 209 358 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00205 561 208 209 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00204 358 211 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00203 211 251 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00202 561 252 211 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00201 561 251 297 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 561 400 190 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00199 190 314 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00198 190 577 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00197 561 184 186 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 186 233 187 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00195 187 185 404 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00194 192 191 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00193 191 271 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00192 561 195 191 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00191 561 323 197 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00190 197 193 195 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00189 195 194 196 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00188 196 233 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00187 561 233 193 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00186 194 323 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00185 561 271 189 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00184 189 314 188 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 561 179 180 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00182 179 577 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00181 561 314 185 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 561 181 182 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 181 314 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00178 183 233 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00177 561 261 183 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00176 561 185 183 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00175 183 400 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00174 561 330 252 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 561 172 118 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00172 118 210 169 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 169 595 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 561 330 114 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 114 289 155 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 171 297 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00167 119 173 172 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 561 171 119 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00165 177 258 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00164 561 330 175 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00163 121 175 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 173 177 121 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 120 330 173 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00160 561 258 120 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 561 155 153 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 561 154 151 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00157 112 153 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00156 113 297 112 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00155 154 192 113 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 115 166 159 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00153 561 330 115 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00152 159 160 157 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00151 561 157 117 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00150 117 160 164 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00149 164 166 116 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00148 160 166 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00147 561 604 166 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00146 116 161 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00145 561 169 161 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00144 330 159 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00143 561 159 330 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 157 164 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00141 111 190 148 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 148 195 111 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 111 151 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 561 130 107 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 107 123 135 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 135 125 106 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 106 136 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 561 136 123 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00133 125 130 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00132 141 595 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00131 561 135 141 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00130 561 183 127 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00129 130 127 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00128 561 128 130 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00127 108 147 138 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00126 561 136 108 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00125 138 145 139 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00124 561 139 109 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00123 109 145 143 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00122 143 147 110 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00121 145 147 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00120 561 604 147 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00119 110 142 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00118 561 141 142 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00117 136 138 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 561 138 136 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 139 143 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00114 561 122 124 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 122 435 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00112 561 252 103 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00111 103 102 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00110 103 297 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00109 105 104 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00108 561 252 105 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 561 103 101 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 101 97 98 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 98 100 99 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 99 104 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 561 104 97 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00102 100 103 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00101 561 96 104 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 96 412 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00099 89 95 88 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00098 561 233 89 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00097 88 94 86 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00096 561 86 87 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00095 87 94 92 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00094 92 95 93 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00093 94 95 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00092 561 604 95 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00091 93 91 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00090 561 90 91 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00089 233 88 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 561 88 233 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 86 92 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00086 90 595 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00085 561 85 90 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00084 561 73 260 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 73 104 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00082 84 233 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00081 561 155 84 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00080 561 251 84 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00079 84 195 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00078 83 84 85 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 85 148 82 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 561 233 81 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00075 81 80 85 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 561 188 83 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 82 233 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 80 184 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00071 561 195 80 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00070 561 76 128 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 78 183 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00068 561 78 79 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 79 78 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 561 128 77 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00065 184 77 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00064 561 136 184 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00063 561 75 74 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 75 136 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00061 70 105 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00060 70 102 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00059 561 251 70 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00058 561 70 71 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 9 51 52 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 561 412 9 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00055 52 50 55 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 561 55 11 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00053 11 50 54 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00052 54 51 10 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00051 50 51 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00050 561 604 51 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00049 10 60 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00048 561 62 60 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 412 52 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 561 52 412 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 55 54 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00044 62 595 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00043 561 98 62 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00042 561 71 12 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 12 64 66 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 66 595 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 561 258 102 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 561 102 13 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 13 251 64 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 6 36 39 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00035 561 251 6 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 39 35 42 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 561 42 8 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 8 35 37 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00031 37 36 7 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00030 35 36 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 561 604 36 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 7 45 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00027 561 66 45 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00026 251 39 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 561 39 251 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 42 37 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 561 79 4 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 4 30 32 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 32 31 5 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 5 76 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 561 76 30 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 31 79 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 561 16 17 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 16 76 561 561 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00015 28 595 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 561 32 28 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 2 19 23 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 561 76 2 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 23 18 21 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 561 21 1 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 1 18 20 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 20 19 3 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 18 19 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 561 604 19 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 3 25 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 561 28 25 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 76 23 561 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 561 23 76 561 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 21 20 561 561 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C603 16 561 1.568e-14
C602 17 561 2.779e-14
C601 18 561 4.869e-14
C600 19 561 5.165e-14
C599 20 561 2.632e-14
C598 21 561 2.005e-14
C596 23 561 2.871e-14
C594 25 561 2.321e-14
C591 28 561 5.402e-14
C589 30 561 2.596e-14
C588 31 561 2.16e-14
C587 32 561 5.214e-14
C586 33 561 7.76e-15
C584 35 561 4.869e-14
C583 36 561 5.165e-14
C582 37 561 2.632e-14
C580 39 561 2.871e-14
C579 40 561 7.33e-15
C578 41 561 7.43e-15
C577 42 561 2.005e-14
C574 45 561 2.321e-14
C569 50 561 4.869e-14
C568 51 561 5.165e-14
C567 52 561 2.871e-14
C565 54 561 2.632e-14
C564 55 561 2.005e-14
C559 60 561 2.321e-14
C557 62 561 5.642e-14
C555 64 561 4.851e-14
C554 65 561 6.05e-15
C553 66 561 8.468e-14
C552 67 561 7.76e-15
C549 70 561 2.455e-14
C548 71 561 6.047e-14
C545 73 561 1.568e-14
C544 74 561 4.603e-14
C543 75 561 1.568e-14
C542 76 561 1.6415e-13
C541 77 561 1.677e-14
C540 78 561 2.552e-14
C539 79 561 6.729e-14
C538 80 561 4.546e-14
C534 84 561 5.656e-14
C533 85 561 6.542e-14
C532 86 561 2.005e-14
C530 88 561 2.871e-14
C528 90 561 6.362e-14
C527 91 561 2.321e-14
C526 92 561 2.632e-14
C524 94 561 4.869e-14
C523 95 561 5.165e-14
C522 96 561 1.568e-14
C521 97 561 2.596e-14
C520 98 561 6.654e-14
C518 100 561 2.16e-14
C516 102 561 1.1547e-13
C515 103 561 6.273e-14
C514 104 561 2.3988e-13
C513 105 561 4.843e-14
C507 111 561 4.11e-15
C495 122 561 1.568e-14
C494 123 561 2.596e-14
C493 124 561 2.899e-14
C492 125 561 2.16e-14
C491 126 561 7.76e-15
C490 127 561 1.677e-14
C489 128 561 8.529e-14
C487 130 561 5.739e-14
C482 135 561 5.454e-14
C481 136 561 1.6028e-13
C479 138 561 2.871e-14
C478 139 561 2.005e-14
C476 141 561 6.122e-14
C475 142 561 2.321e-14
C474 143 561 2.632e-14
C472 145 561 4.869e-14
C470 147 561 5.165e-14
C469 148 561 5.327e-14
C466 151 561 5.535e-14
C464 153 561 4.599e-14
C463 154 561 2.605e-14
C462 155 561 8.727e-14
C461 156 561 7.76e-15
C460 157 561 2.005e-14
C458 159 561 2.871e-14
C457 160 561 4.869e-14
C456 161 561 2.321e-14
C453 164 561 2.632e-14
C451 166 561 5.165e-14
C448 169 561 5.348e-14
C447 170 561 6.05e-15
C446 171 561 1.662e-14
C445 172 561 4.581e-14
C444 173 561 5.7e-14
C443 174 561 9.7e-15
C442 175 561 2.596e-14
C440 177 561 2.16e-14
C437 179 561 1.568e-14
C436 180 561 4.003e-14
C435 181 561 1.568e-14
C434 182 561 3.667e-14
C433 183 561 1.125e-13
C432 184 561 1.0867e-13
C431 185 561 8.23e-14
C428 188 561 6.264e-14
C426 190 561 5.347e-14
C425 191 561 1.8635e-14
C424 192 561 5.231e-14
C423 193 561 2.596e-14
C422 194 561 2.16e-14
C421 195 561 1.7436e-13
C418 198 561 2.871e-14
C416 200 561 2.005e-14
C414 202 561 2.632e-14
C412 204 561 2.321e-14
C411 205 561 4.869e-14
C410 206 561 5.165e-14
C409 207 561 1.568e-14
C408 208 561 5.053e-14
C407 209 561 1.8635e-14
C406 210 561 6.461e-14
C405 211 561 1.8635e-14
C393 222 561 1.568e-14
C392 223 561 1.568e-14
C391 224 561 2.371e-14
C390 225 561 3.547e-14
C389 226 561 1.568e-14
C388 227 561 1.568e-14
C387 228 561 4.507e-14
C386 229 561 1.8635e-14
C385 230 561 9.7e-15
C384 231 561 2.596e-14
C383 232 561 6.369e-14
C382 233 561 4.12101e-13
C381 234 561 2.16e-14
C380 235 561 2.005e-14
C379 236 561 2.632e-14
C376 239 561 2.871e-14
C375 240 561 2.321e-14
C373 242 561 4.869e-14
C372 243 561 5.165e-14
C371 244 561 1.662e-14
C370 245 561 5.211e-14
C369 246 561 5.468e-14
C368 247 561 6.05e-15
C367 248 561 4.581e-14
C366 249 561 1.8635e-14
C365 250 561 9.438e-14
C364 251 561 4.6844e-13
C363 252 561 1.5885e-13
C359 256 561 5.247e-14
C358 257 561 1.677e-14
C357 258 561 1.2774e-13
C355 260 561 7.867e-14
C354 261 561 8.562e-14
C347 268 561 5.01e-14
C344 271 561 1.4509e-13
C340 275 561 6.05e-15
C339 276 561 6.428e-14
C336 279 561 1.662e-14
C334 281 561 9.7e-15
C332 283 561 6.06e-14
C329 286 561 5.246e-14
C326 289 561 1.5659e-13
C321 293 561 9.7e-15
C318 296 561 8.148e-14
C317 297 561 3.1656e-13
C316 298 561 2.306e-14
C314 300 561 2.605e-14
C310 304 561 1.8635e-14
C309 305 561 1.3755e-13
C308 306 561 4.11e-15
C307 307 561 4.581e-14
C306 308 561 5.625e-14
C303 311 561 2.596e-14
C302 312 561 2.16e-14
C300 314 561 3.3082e-13
C299 315 561 5.817e-14
C296 318 561 2.306e-14
C295 319 561 1.568e-14
C294 320 561 2.596e-14
C293 321 561 2.16e-14
C292 322 561 6.133e-14
C291 323 561 4.3378e-13
C289 324 561 2.659e-14
C288 325 561 1.568e-14
C287 326 561 5.925e-14
C284 329 561 5.226e-14
C283 330 561 3.6787e-13
C282 331 561 6.026e-14
C281 332 561 9.155e-14
C279 334 561 1.677e-14
C278 335 561 7.375e-14
C277 336 561 1.853e-14
C275 338 561 2.8915e-13
C273 340 561 2.871e-14
C272 341 561 2.005e-14
C270 343 561 2.632e-14
C269 344 561 7.038e-14
C268 345 561 2.321e-14
C266 347 561 4.869e-14
C265 348 561 5.165e-14
C264 349 561 1.1506e-13
C262 351 561 1.677e-14
C261 352 561 6.058e-14
C260 353 561 5.008e-14
C259 354 561 9.779e-14
C257 356 561 1.568e-14
C256 357 561 8.311e-14
C255 358 561 1.0938e-13
C252 361 561 1.2764e-13
C251 362 561 1.1617e-13
C250 363 561 6.835e-14
C242 371 561 7.185e-14
C237 376 561 1.7866e-13
C229 383 561 7.76e-15
C228 384 561 1.2819e-13
C227 385 561 2.306e-14
C224 388 561 4.779e-14
C222 390 561 1.1695e-13
C221 391 561 1.8635e-14
C217 395 561 6.75e-14
C216 396 561 5.938e-14
C215 397 561 4.828e-14
C214 398 561 1.8635e-14
C212 400 561 1.7261e-13
C211 401 561 2.455e-14
C208 404 561 1.527e-13
C207 405 561 1.568e-14
C206 406 561 1.568e-14
C205 407 561 1.0497e-13
C204 408 561 9.883e-14
C200 412 561 2.0081e-13
C199 413 561 2.871e-14
C197 415 561 4.869e-14
C196 416 561 2.632e-14
C194 418 561 2.005e-14
C193 419 561 2.321e-14
C192 420 561 5.642e-14
C191 421 561 5.165e-14
C189 423 561 2.596e-14
C188 424 561 2.16e-14
C187 425 561 3.4951e-13
C186 426 561 5.454e-14
C182 429 561 1.0512e-13
C181 430 561 1.568e-14
C180 431 561 2.596e-14
C179 432 561 6.009e-14
C178 433 561 2.16e-14
C177 434 561 9.7e-15
C176 435 561 2.4507e-13
C175 436 561 2.871e-14
C173 438 561 2.005e-14
C171 440 561 2.632e-14
C169 442 561 7.26e-14
C168 443 561 2.321e-14
C167 444 561 4.869e-14
C166 445 561 5.165e-14
C165 446 561 1.662e-14
C164 447 561 4.941e-14
C163 448 561 5.309e-14
C162 449 561 5.674e-14
C161 450 561 5.708e-14
C160 451 561 5.361e-14
C159 452 561 6.05e-15
C158 453 561 1.662e-14
C156 455 561 2.871e-14
C155 456 561 2.005e-14
C153 458 561 2.632e-14
C152 459 561 2.321e-14
C150 461 561 4.869e-14
C149 462 561 1.1621e-13
C148 463 561 5.165e-14
C147 464 561 1.568e-14
C146 465 561 1.8635e-14
C145 466 561 9.849e-14
C143 468 561 2.455e-14
C141 470 561 5.447e-14
C140 471 561 6.908e-14
C139 472 561 6.05e-15
C138 473 561 4.421e-14
C136 475 561 1.8635e-14
C133 478 561 2.455e-14
C132 479 561 6.76e-14
C128 483 561 1.2966e-13
C123 488 561 9.7e-15
C122 489 561 6.05e-15
C120 491 561 6.05e-15
C119 492 561 9.7e-15
C118 493 561 6.05e-15
C113 497 561 3.139e-14
C112 498 561 1.568e-14
C111 499 561 3.187e-14
C110 500 561 1.568e-14
C108 502 561 2.005e-14
C107 503 561 2.871e-14
C105 505 561 2.321e-14
C103 507 561 2.632e-14
C100 510 561 4.869e-14
C99 511 561 5.165e-14
C97 513 561 1.2877e-13
C96 514 561 1.6417e-13
C95 515 561 1.8635e-14
C93 517 561 3.9674e-13
C92 518 561 2.596e-14
C89 521 561 5.1e-14
C88 522 561 1.662e-14
C86 524 561 2.16e-14
C83 527 561 7.988e-14
C80 530 561 2.0454e-13
C79 531 561 1.8635e-14
C78 532 561 4.421e-14
C77 533 561 8.117e-14
C76 534 561 6.257e-14
C74 536 561 1.767e-14
C73 537 561 5.087e-14
C72 538 561 3.1843e-13
C70 540 561 2.596e-14
C68 542 561 5.1e-14
C67 543 561 1.662e-14
C65 545 561 2.16e-14
C64 546 561 4.941e-14
C59 551 561 2.632e-14
C58 552 561 2.871e-14
C57 553 561 2.005e-14
C55 555 561 6.068e-14
C53 557 561 2.321e-14
C52 558 561 4.869e-14
C51 559 561 5.165e-14
C49 561 561 6.78197e-12
C48 562 561 1.568e-14
C47 563 561 2.659e-14
C46 564 561 1.2576e-13
C45 565 561 1.568e-14
C44 566 561 2.596e-14
C43 567 561 6.249e-14
C42 568 561 2.16e-14
C41 569 561 9.7e-15
C40 570 561 5.34e-14
C39 571 561 1.6343e-13
C38 572 561 1.662e-14
C37 573 561 5.141e-14
C36 574 561 5.181e-14
C35 575 561 6.05e-15
C33 577 561 3.4558e-13
C32 578 561 2.871e-14
C31 579 561 2.005e-14
C29 581 561 2.632e-14
C28 582 561 6.308e-14
C27 583 561 2.321e-14
C25 585 561 4.869e-14
C24 586 561 5.165e-14
C23 587 561 1.568e-14
C22 588 561 1.1035e-13
C21 589 561 2.4917e-13
C20 590 561 1.8635e-14
C18 592 561 6.941e-14
C17 593 561 3.7268e-13
C16 594 561 3.7629e-13
C15 595 561 8.65419e-13
C12 598 561 6.0004e-13
C11 599 561 2.871e-14
C10 600 561 2.005e-14
C8 602 561 2.632e-14
C7 603 561 6.482e-14
C6 604 561 8.65549e-13
C4 606 561 2.321e-14
C3 607 561 4.869e-14
C2 608 561 7.1205e-12
C1 609 561 5.165e-14
.ends act4_cougar

