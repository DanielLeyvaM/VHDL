* Spice description of sum4b_cougar
* Spice driver version -1208856924
* Date ( dd/mm/yyyy hh:mm:ss ):  9/10/2020 at 20:36:57

* INTERF a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] ci co so[0] so[1] so[2] 
* INTERF so[3] vdd vss 


.subckt sum4b_cougar a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] ci co so[0] so[1] so[2] so[3] vdd vss 
Mtr_00154 acarreo0 sig4 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00153 sig2 a[0] sig3 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00152 sig2 b[0] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00151 vdd a[0] sig2 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00150 sig3 b[0] sig4 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00149 sig4 cix sig2 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00148 sig13 b[0] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 vdd a[0] sig10 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 x0.xr2_x1_sig sig13 sig11 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00145 sig11 a[0] vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00144 sig11 sig10 x0.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00143 vdd b[0] sig11 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00142 sig19 cix vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 vdd x0.xr2_x1_sig sig16 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 so[0] sig19 sig17 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00139 sig17 x0.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00138 sig17 sig16 so[0] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00137 vdd cix sig17 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00136 sig36 b[1] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 vdd a[1] sig31 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 x1.xr2_x1_sig sig36 sig47 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00133 sig47 a[1] vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00132 sig47 sig31 x1.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00131 vdd b[1] sig47 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00130 acarreo1 sig25 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00129 sig45 a[1] sig46 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00128 sig45 b[1] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00127 vdd a[1] sig45 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00126 sig46 b[1] sig25 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00125 sig25 acarreo0 sig45 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00124 vdd ci sig22 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00123 vdd sig22 cix vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00122 cix sig22 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00121 vdd sig22 cix vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00120 cix sig22 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00119 sig43 acarreo0 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 vdd x1.xr2_x1_sig sig39 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 so[1] sig43 sig48 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00116 sig48 x1.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00115 sig48 sig39 so[1] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00114 vdd acarreo0 sig48 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00113 sig52 b[2] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 vdd a[2] sig49 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 x2.xr2_x1_sig sig52 sig51 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00110 sig51 a[2] vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00109 sig51 sig49 x2.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00108 vdd b[2] sig51 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00107 sig57 acarreo1 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 vdd x2.xr2_x1_sig sig54 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 so[2] sig57 sig55 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00104 sig55 x2.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00103 sig55 sig54 so[2] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00102 vdd acarreo1 sig55 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00101 sig62 b[3] vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 vdd a[3] sig58 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 x3.xr2_x1_sig sig62 sig60 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00098 sig60 a[3] vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00097 sig60 sig58 x3.xr2_x1_sig vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00096 vdd b[3] sig60 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00095 sig66 acarreo2 vdd vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 vdd x3.xr2_x1_sig sig64 vdd tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 so[3] sig66 sig63 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00092 sig63 x3.xr2_x1_sig vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00091 sig63 sig64 so[3] vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00090 vdd acarreo2 sig63 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00089 acarreo2 sig72 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00088 sig81 a[2] sig83 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00087 sig81 b[2] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00086 vdd a[2] sig81 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00085 sig83 b[2] sig72 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00084 sig72 acarreo1 sig81 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00083 co sig77 vdd vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00082 sig84 a[3] sig87 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00081 sig84 b[3] vdd vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00080 vdd a[3] sig84 vdd tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00079 sig87 b[3] sig77 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00078 sig77 acarreo2 sig84 vdd tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00077 vss sig4 acarreo0 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 vss b[0] sig20 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00075 sig20 a[0] vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00074 sig4 b[0] sig23 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00073 sig23 a[0] vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00072 sig20 cix sig4 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00071 sig10 a[0] vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00070 vss b[0] sig13 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 sig32 sig13 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 x0.xr2_x1_sig sig10 sig32 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 sig29 b[0] x0.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 vss a[0] sig29 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 sig16 x0.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00064 vss cix sig19 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00063 sig37 sig19 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 so[0] sig16 sig37 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 sig38 cix so[0] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 vss x0.xr2_x1_sig sig38 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 sig31 a[1] vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00058 vss b[1] sig36 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00057 sig33 sig36 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 x1.xr2_x1_sig sig31 sig33 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 sig34 b[1] x1.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 vss a[1] sig34 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 vss sig25 acarreo1 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 vss b[1] sig27 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00051 sig27 a[1] vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00050 sig25 b[1] sig26 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00049 sig26 a[1] vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00048 sig27 acarreo0 sig25 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00047 sig22 ci vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 cix sig22 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 vss sig22 cix vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 vss sig22 cix vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 cix sig22 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 sig39 x1.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00041 vss acarreo0 sig43 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00040 sig42 sig43 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 so[1] sig39 sig42 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 sig40 acarreo0 so[1] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 vss x1.xr2_x1_sig sig40 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 sig49 a[2] vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00035 vss b[2] sig52 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 sig68 sig52 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 x2.xr2_x1_sig sig49 sig68 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 sig70 b[2] x2.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 vss a[2] sig70 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 sig54 x2.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 vss acarreo1 sig57 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 sig73 sig57 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 so[2] sig54 sig73 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 sig71 acarreo1 so[2] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 vss x2.xr2_x1_sig sig71 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 sig58 a[3] vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 vss b[3] sig62 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 sig74 sig62 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 x3.xr2_x1_sig sig58 sig74 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 sig75 b[3] x3.xr2_x1_sig vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 vss a[3] sig75 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 sig64 x3.xr2_x1_sig vss vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 vss acarreo2 sig66 vss tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 sig78 sig66 vss vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 so[3] sig64 sig78 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 sig76 acarreo2 so[3] vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 vss x3.xr2_x1_sig sig76 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 vss sig72 acarreo2 vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 vss b[2] sig79 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00010 sig79 a[2] vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00009 sig72 b[2] sig80 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00008 sig80 a[2] vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00007 sig79 acarreo1 sig72 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00006 vss sig77 co vss tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 vss b[3] sig85 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00004 sig85 a[3] vss vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00003 sig77 b[3] sig86 vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00002 sig86 a[3] vss vss tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00001 sig85 acarreo2 sig77 vss tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
C88 co vss 2.816e-14
C85 sig85 vss 4.11e-15
C84 sig84 vss 8.58e-15
C81 sig81 vss 8.58e-15
C79 sig79 vss 4.11e-15
C77 sig77 vss 2.299e-14
C72 sig72 vss 2.299e-14
C67 acarreo2 vss 1.1581e-13
C66 sig66 vss 2.596e-14
C65 so[3] vss 3.889e-14
C64 sig64 vss 2.16e-14
C63 sig63 vss 9.7e-15
C62 sig62 vss 2.596e-14
C61 a[3] vss 1.0814e-13
C60 sig60 vss 9.7e-15
C59 x3.xr2_x1_sig vss 5.751e-14
C58 sig58 vss 2.16e-14
C57 sig57 vss 2.596e-14
C56 so[2] vss 5.281e-14
C55 sig55 vss 9.7e-15
C54 sig54 vss 2.16e-14
C53 a[2] vss 8.534e-14
C52 sig52 vss 2.596e-14
C51 sig51 vss 9.7e-15
C50 x2.xr2_x1_sig vss 5.751e-14
C49 sig49 vss 2.16e-14
C48 sig48 vss 9.7e-15
C47 sig47 vss 9.7e-15
C45 sig45 vss 8.58e-15
C43 sig43 vss 2.596e-14
C41 so[1] vss 3.409e-14
C39 sig39 vss 2.16e-14
C36 sig36 vss 2.596e-14
C35 x1.xr2_x1_sig vss 5.751e-14
C31 sig31 vss 2.16e-14
C30 acarreo1 vss 1.0909e-13
C28 a[1] vss 8.862e-14
C27 sig27 vss 4.11e-15
C25 sig25 vss 2.299e-14
C24 ci vss 6.429e-14
C22 sig22 vss 4.103e-14
C21 vss vss 8.34002e-13
C20 sig20 vss 4.11e-15
C19 sig19 vss 2.596e-14
C18 so[0] vss 3.649e-14
C17 sig17 vss 9.7e-15
C16 sig16 vss 2.16e-14
C15 b[3] vss 1.3016e-13
C14 b[2] vss 1.3728e-13
C13 sig13 vss 2.596e-14
C12 x0.xr2_x1_sig vss 5.991e-14
C11 sig11 vss 9.7e-15
C10 sig10 vss 2.16e-14
C9 b[1] vss 1.032e-13
C8 acarreo0 vss 1.1053e-13
C7 a[0] vss 8.262e-14
C6 b[0] vss 9.552e-14
C5 cix vss 1.2765e-13
C4 sig4 vss 2.299e-14
C2 sig2 vss 8.58e-15
C1 vdd vss 8.44081e-13
.ends sum4b_cougar

